`timescale 1ns / 1ps
module bmpsimplifyinput_rom (
    input wire clk,
    input wire [7:0] row,
    input wire [9:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 640 + col) >= 0 && (row * 640 + col) <= 12180) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 12181 && (row * 640 + col) <= 12307) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 12308 && (row * 640 + col) <= 12336) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 12337 && (row * 640 + col) <= 12465) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 12466 && (row * 640 + col) <= 12728) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 12729 && (row * 640 + col) <= 12735) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 12736 && (row * 640 + col) <= 12817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 12818 && (row * 640 + col) <= 12950) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 12951 && (row * 640 + col) <= 12974) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 12975 && (row * 640 + col) <= 13108) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 13109 && (row * 640 + col) <= 13365) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 13366 && (row * 640 + col) <= 13382) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 13383 && (row * 640 + col) <= 13455) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 13456 && (row * 640 + col) <= 13592) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 13593 && (row * 640 + col) <= 13612) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 13613 && (row * 640 + col) <= 13750) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 13751 && (row * 640 + col) <= 14004) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14005 && (row * 640 + col) <= 14025) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 14026 && (row * 640 + col) <= 14093) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14094 && (row * 640 + col) <= 14233) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 14234 && (row * 640 + col) <= 14251) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14252 && (row * 640 + col) <= 14391) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 14392 && (row * 640 + col) <= 14643) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14644 && (row * 640 + col) <= 14668) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 14669 && (row * 640 + col) <= 14732) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14733 && (row * 640 + col) <= 14874) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 14875 && (row * 640 + col) <= 14890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14891 && (row * 640 + col) <= 15032) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 15033 && (row * 640 + col) <= 15282) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 15283 && (row * 640 + col) <= 15310) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 15311 && (row * 640 + col) <= 15371) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 15372 && (row * 640 + col) <= 15515) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 15516 && (row * 640 + col) <= 15529) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 15530 && (row * 640 + col) <= 15673) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 15674 && (row * 640 + col) <= 15922) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 15923 && (row * 640 + col) <= 15952) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 15953 && (row * 640 + col) <= 16011) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16012 && (row * 640 + col) <= 16156) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 16157 && (row * 640 + col) <= 16168) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16169 && (row * 640 + col) <= 16314) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 16315 && (row * 640 + col) <= 16562) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16563 && (row * 640 + col) <= 16568) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 16569 && (row * 640 + col) <= 16578) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16579 && (row * 640 + col) <= 16595) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 16596 && (row * 640 + col) <= 16650) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16651 && (row * 640 + col) <= 16797) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 16798 && (row * 640 + col) <= 16808) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16809 && (row * 640 + col) <= 16955) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 16956 && (row * 640 + col) <= 17202) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17203 && (row * 640 + col) <= 17207) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 17208 && (row * 640 + col) <= 17222) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17223 && (row * 640 + col) <= 17236) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 17237 && (row * 640 + col) <= 17289) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17290 && (row * 640 + col) <= 17300) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17301 && (row * 640 + col) <= 17428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17429 && (row * 640 + col) <= 17437) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17438 && (row * 640 + col) <= 17447) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17448 && (row * 640 + col) <= 17457) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17458 && (row * 640 + col) <= 17585) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17586 && (row * 640 + col) <= 17595) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17596 && (row * 640 + col) <= 17842) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17843 && (row * 640 + col) <= 17847) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 17848 && (row * 640 + col) <= 17866) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17867 && (row * 640 + col) <= 17878) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 17879 && (row * 640 + col) <= 17929) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17930 && (row * 640 + col) <= 17938) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17939 && (row * 640 + col) <= 18069) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18070 && (row * 640 + col) <= 18078) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18079 && (row * 640 + col) <= 18087) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18088 && (row * 640 + col) <= 18095) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18096 && (row * 640 + col) <= 18227) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18228 && (row * 640 + col) <= 18236) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18237 && (row * 640 + col) <= 18301) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18302 && (row * 640 + col) <= 18313) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18314 && (row * 640 + col) <= 18482) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18483 && (row * 640 + col) <= 18488) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 18489 && (row * 640 + col) <= 18508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18509 && (row * 640 + col) <= 18520) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 18521 && (row * 640 + col) <= 18569) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18570 && (row * 640 + col) <= 18577) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18578 && (row * 640 + col) <= 18710) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18711 && (row * 640 + col) <= 18718) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18719 && (row * 640 + col) <= 18726) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18727 && (row * 640 + col) <= 18734) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18735 && (row * 640 + col) <= 18868) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18869 && (row * 640 + col) <= 18876) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18877 && (row * 640 + col) <= 18939) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18940 && (row * 640 + col) <= 18955) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18956 && (row * 640 + col) <= 19122) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19123 && (row * 640 + col) <= 19130) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 19131 && (row * 640 + col) <= 19150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19151 && (row * 640 + col) <= 19161) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 19162 && (row * 640 + col) <= 19208) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19209 && (row * 640 + col) <= 19216) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19217 && (row * 640 + col) <= 19351) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19352 && (row * 640 + col) <= 19358) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19359 && (row * 640 + col) <= 19366) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19367 && (row * 640 + col) <= 19374) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19375 && (row * 640 + col) <= 19508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19509 && (row * 640 + col) <= 19516) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19517 && (row * 640 + col) <= 19577) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19578 && (row * 640 + col) <= 19598) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19599 && (row * 640 + col) <= 19763) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19764 && (row * 640 + col) <= 19773) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 19774 && (row * 640 + col) <= 19792) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19793 && (row * 640 + col) <= 19802) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 19803 && (row * 640 + col) <= 19848) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19849 && (row * 640 + col) <= 19856) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19857 && (row * 640 + col) <= 19991) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19992 && (row * 640 + col) <= 19999) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20000 && (row * 640 + col) <= 20006) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20007 && (row * 640 + col) <= 20013) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20014 && (row * 640 + col) <= 20149) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20150 && (row * 640 + col) <= 20156) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20157 && (row * 640 + col) <= 20215) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20216 && (row * 640 + col) <= 20239) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20240 && (row * 640 + col) <= 20403) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20404 && (row * 640 + col) <= 20415) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 20416 && (row * 640 + col) <= 20434) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20435 && (row * 640 + col) <= 20444) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 20445 && (row * 640 + col) <= 20488) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20489 && (row * 640 + col) <= 20495) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20496 && (row * 640 + col) <= 20631) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20632 && (row * 640 + col) <= 20639) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20640 && (row * 640 + col) <= 20646) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20647 && (row * 640 + col) <= 20653) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20654 && (row * 640 + col) <= 20789) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20790 && (row * 640 + col) <= 20797) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20798 && (row * 640 + col) <= 20854) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20855 && (row * 640 + col) <= 20880) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20881 && (row * 640 + col) <= 21044) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21045 && (row * 640 + col) <= 21056) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 21057 && (row * 640 + col) <= 21075) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21076 && (row * 640 + col) <= 21085) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 21086 && (row * 640 + col) <= 21128) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21129 && (row * 640 + col) <= 21135) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21136 && (row * 640 + col) <= 21271) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21272 && (row * 640 + col) <= 21279) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21280 && (row * 640 + col) <= 21286) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21287 && (row * 640 + col) <= 21293) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21294 && (row * 640 + col) <= 21429) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21430 && (row * 640 + col) <= 21437) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21438 && (row * 640 + col) <= 21493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21494 && (row * 640 + col) <= 21522) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21523 && (row * 640 + col) <= 21686) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21687 && (row * 640 + col) <= 21698) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 21699 && (row * 640 + col) <= 21717) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21718 && (row * 640 + col) <= 21726) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 21727 && (row * 640 + col) <= 21768) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21769 && (row * 640 + col) <= 21775) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21776 && (row * 640 + col) <= 21911) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21912 && (row * 640 + col) <= 21919) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21920 && (row * 640 + col) <= 21926) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21927 && (row * 640 + col) <= 21933) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21934 && (row * 640 + col) <= 22069) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22070 && (row * 640 + col) <= 22077) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22078 && (row * 640 + col) <= 22132) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22133 && (row * 640 + col) <= 22163) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22164 && (row * 640 + col) <= 22328) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22329 && (row * 640 + col) <= 22340) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 22341 && (row * 640 + col) <= 22358) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22359 && (row * 640 + col) <= 22367) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 22368 && (row * 640 + col) <= 22408) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22409 && (row * 640 + col) <= 22415) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22416 && (row * 640 + col) <= 22551) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22552 && (row * 640 + col) <= 22559) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22560 && (row * 640 + col) <= 22566) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22567 && (row * 640 + col) <= 22573) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22574 && (row * 640 + col) <= 22709) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22710 && (row * 640 + col) <= 22716) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22717 && (row * 640 + col) <= 22771) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22772 && (row * 640 + col) <= 22804) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22805 && (row * 640 + col) <= 22970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22971 && (row * 640 + col) <= 22982) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 22983 && (row * 640 + col) <= 23000) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23001 && (row * 640 + col) <= 23008) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 23009 && (row * 640 + col) <= 23048) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23049 && (row * 640 + col) <= 23056) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23057 && (row * 640 + col) <= 23191) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23192 && (row * 640 + col) <= 23198) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23199 && (row * 640 + col) <= 23206) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23207 && (row * 640 + col) <= 23214) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23215 && (row * 640 + col) <= 23348) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23349 && (row * 640 + col) <= 23356) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23357 && (row * 640 + col) <= 23410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23411 && (row * 640 + col) <= 23423) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23424 && (row * 640 + col) <= 23432) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23433 && (row * 640 + col) <= 23444) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23445 && (row * 640 + col) <= 23612) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23613 && (row * 640 + col) <= 23623) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 23624 && (row * 640 + col) <= 23641) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23642 && (row * 640 + col) <= 23649) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 23650 && (row * 640 + col) <= 23688) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23689 && (row * 640 + col) <= 23696) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23697 && (row * 640 + col) <= 23830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23831 && (row * 640 + col) <= 23838) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23839 && (row * 640 + col) <= 23846) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23847 && (row * 640 + col) <= 23854) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23855 && (row * 640 + col) <= 23988) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23989 && (row * 640 + col) <= 23996) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23997 && (row * 640 + col) <= 24049) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24050 && (row * 640 + col) <= 24061) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24062 && (row * 640 + col) <= 24074) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24075 && (row * 640 + col) <= 24085) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24086 && (row * 640 + col) <= 24254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24255 && (row * 640 + col) <= 24265) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 24266 && (row * 640 + col) <= 24282) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24283 && (row * 640 + col) <= 24290) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 24291 && (row * 640 + col) <= 24329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24330 && (row * 640 + col) <= 24337) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24338 && (row * 640 + col) <= 24470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24471 && (row * 640 + col) <= 24478) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24479 && (row * 640 + col) <= 24486) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24487 && (row * 640 + col) <= 24495) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24496 && (row * 640 + col) <= 24627) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24628 && (row * 640 + col) <= 24636) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24637 && (row * 640 + col) <= 24689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24690 && (row * 640 + col) <= 24699) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24700 && (row * 640 + col) <= 24716) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24717 && (row * 640 + col) <= 24726) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24727 && (row * 640 + col) <= 24896) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24897 && (row * 640 + col) <= 24906) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 24907 && (row * 640 + col) <= 24923) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24924 && (row * 640 + col) <= 24931) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 24932 && (row * 640 + col) <= 24969) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24970 && (row * 640 + col) <= 24978) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24979 && (row * 640 + col) <= 25108) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25109 && (row * 640 + col) <= 25118) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25119 && (row * 640 + col) <= 25127) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25128 && (row * 640 + col) <= 25136) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25137 && (row * 640 + col) <= 25266) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25267 && (row * 640 + col) <= 25275) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25276 && (row * 640 + col) <= 25328) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25329 && (row * 640 + col) <= 25338) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25339 && (row * 640 + col) <= 25357) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25358 && (row * 640 + col) <= 25366) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25367 && (row * 640 + col) <= 25474) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25475 && (row * 640 + col) <= 25491) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25492 && (row * 640 + col) <= 25537) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25538 && (row * 640 + col) <= 25548) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 25549 && (row * 640 + col) <= 25564) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25565 && (row * 640 + col) <= 25572) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 25573 && (row * 640 + col) <= 25610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25611 && (row * 640 + col) <= 25619) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25620 && (row * 640 + col) <= 25746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25747 && (row * 640 + col) <= 25757) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25758 && (row * 640 + col) <= 25767) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25768 && (row * 640 + col) <= 25778) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25779 && (row * 640 + col) <= 25904) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25905 && (row * 640 + col) <= 25915) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25916 && (row * 640 + col) <= 25968) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25969 && (row * 640 + col) <= 25977) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25978 && (row * 640 + col) <= 25998) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25999 && (row * 640 + col) <= 26007) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26008 && (row * 640 + col) <= 26107) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26108 && (row * 640 + col) <= 26136) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26137 && (row * 640 + col) <= 26179) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26180 && (row * 640 + col) <= 26189) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 26190 && (row * 640 + col) <= 26205) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26206 && (row * 640 + col) <= 26213) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 26214 && (row * 640 + col) <= 26250) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26251 && (row * 640 + col) <= 26396) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26397 && (row * 640 + col) <= 26408) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26409 && (row * 640 + col) <= 26554) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26555 && (row * 640 + col) <= 26607) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26608 && (row * 640 + col) <= 26616) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26617 && (row * 640 + col) <= 26638) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26639 && (row * 640 + col) <= 26647) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26648 && (row * 640 + col) <= 26741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26742 && (row * 640 + col) <= 26780) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26781 && (row * 640 + col) <= 26821) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26822 && (row * 640 + col) <= 26831) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 26832 && (row * 640 + col) <= 26846) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26847 && (row * 640 + col) <= 26854) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 26855 && (row * 640 + col) <= 26891) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26892 && (row * 640 + col) <= 27036) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27037 && (row * 640 + col) <= 27048) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27049 && (row * 640 + col) <= 27194) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27195 && (row * 640 + col) <= 27247) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27248 && (row * 640 + col) <= 27256) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27257 && (row * 640 + col) <= 27279) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27280 && (row * 640 + col) <= 27287) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27288 && (row * 640 + col) <= 27378) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27379 && (row * 640 + col) <= 27422) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27423 && (row * 640 + col) <= 27462) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27463 && (row * 640 + col) <= 27472) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 27473 && (row * 640 + col) <= 27487) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27488 && (row * 640 + col) <= 27494) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 27495 && (row * 640 + col) <= 27532) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27533 && (row * 640 + col) <= 27675) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27676 && (row * 640 + col) <= 27689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27690 && (row * 640 + col) <= 27833) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27834 && (row * 640 + col) <= 27887) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27888 && (row * 640 + col) <= 27895) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27896 && (row * 640 + col) <= 27920) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27921 && (row * 640 + col) <= 27928) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27929 && (row * 640 + col) <= 28015) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28016 && (row * 640 + col) <= 28065) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28066 && (row * 640 + col) <= 28104) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28105 && (row * 640 + col) <= 28113) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 28114 && (row * 640 + col) <= 28128) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28129 && (row * 640 + col) <= 28135) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 28136 && (row * 640 + col) <= 28173) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28174 && (row * 640 + col) <= 28314) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28315 && (row * 640 + col) <= 28330) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28331 && (row * 640 + col) <= 28472) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28473 && (row * 640 + col) <= 28526) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28527 && (row * 640 + col) <= 28535) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28536 && (row * 640 + col) <= 28560) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28561 && (row * 640 + col) <= 28568) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28569 && (row * 640 + col) <= 28652) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28653 && (row * 640 + col) <= 28707) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28708 && (row * 640 + col) <= 28745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28746 && (row * 640 + col) <= 28755) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 28756 && (row * 640 + col) <= 28769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28770 && (row * 640 + col) <= 28776) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 28777 && (row * 640 + col) <= 28814) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28815 && (row * 640 + col) <= 28953) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28954 && (row * 640 + col) <= 28971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28972 && (row * 640 + col) <= 29111) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29112 && (row * 640 + col) <= 29166) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29167 && (row * 640 + col) <= 29174) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29175 && (row * 640 + col) <= 29200) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29201 && (row * 640 + col) <= 29208) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29209 && (row * 640 + col) <= 29290) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29291 && (row * 640 + col) <= 29348) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29349 && (row * 640 + col) <= 29387) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29388 && (row * 640 + col) <= 29396) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 29397 && (row * 640 + col) <= 29410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29411 && (row * 640 + col) <= 29416) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 29417 && (row * 640 + col) <= 29455) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29456 && (row * 640 + col) <= 29591) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29592 && (row * 640 + col) <= 29613) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29614 && (row * 640 + col) <= 29749) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29750 && (row * 640 + col) <= 29806) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29807 && (row * 640 + col) <= 29814) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29815 && (row * 640 + col) <= 29840) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29841 && (row * 640 + col) <= 29848) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29849 && (row * 640 + col) <= 29927) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29928 && (row * 640 + col) <= 29990) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29991 && (row * 640 + col) <= 30028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30029 && (row * 640 + col) <= 30037) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 30038 && (row * 640 + col) <= 30050) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30051 && (row * 640 + col) <= 30057) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 30058 && (row * 640 + col) <= 30097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30098 && (row * 640 + col) <= 30229) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 30230 && (row * 640 + col) <= 30255) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30256 && (row * 640 + col) <= 30387) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 30388 && (row * 640 + col) <= 30446) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30447 && (row * 640 + col) <= 30454) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 30455 && (row * 640 + col) <= 30480) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30481 && (row * 640 + col) <= 30488) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 30489 && (row * 640 + col) <= 30566) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30567 && (row * 640 + col) <= 30631) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 30632 && (row * 640 + col) <= 30669) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30670 && (row * 640 + col) <= 30678) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 30679 && (row * 640 + col) <= 30691) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30692 && (row * 640 + col) <= 30698) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 30699 && (row * 640 + col) <= 30899) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30900 && (row * 640 + col) <= 31023) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31024 && (row * 640 + col) <= 31086) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31087 && (row * 640 + col) <= 31094) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31095 && (row * 640 + col) <= 31120) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31121 && (row * 640 + col) <= 31128) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31129 && (row * 640 + col) <= 31204) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31205 && (row * 640 + col) <= 31232) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31233 && (row * 640 + col) <= 31252) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31253 && (row * 640 + col) <= 31272) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31273 && (row * 640 + col) <= 31311) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31312 && (row * 640 + col) <= 31319) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 31320 && (row * 640 + col) <= 31332) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31333 && (row * 640 + col) <= 31338) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 31339 && (row * 640 + col) <= 31726) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31727 && (row * 640 + col) <= 31734) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31735 && (row * 640 + col) <= 31760) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31761 && (row * 640 + col) <= 31768) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31769 && (row * 640 + col) <= 31842) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31843 && (row * 640 + col) <= 31865) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31866 && (row * 640 + col) <= 31897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31898 && (row * 640 + col) <= 31913) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31914 && (row * 640 + col) <= 31952) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31953 && (row * 640 + col) <= 31961) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 31962 && (row * 640 + col) <= 31972) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31973 && (row * 640 + col) <= 31979) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 31980 && (row * 640 + col) <= 32366) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32367 && (row * 640 + col) <= 32374) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 32375 && (row * 640 + col) <= 32400) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32401 && (row * 640 + col) <= 32408) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 32409 && (row * 640 + col) <= 32481) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32482 && (row * 640 + col) <= 32502) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 32503 && (row * 640 + col) <= 32539) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32540 && (row * 640 + col) <= 32553) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 32554 && (row * 640 + col) <= 32593) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32594 && (row * 640 + col) <= 32602) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 32603 && (row * 640 + col) <= 32613) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32614 && (row * 640 + col) <= 32619) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 32620 && (row * 640 + col) <= 33006) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33007 && (row * 640 + col) <= 33014) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33015 && (row * 640 + col) <= 33040) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33041 && (row * 640 + col) <= 33048) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33049 && (row * 640 + col) <= 33119) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33120 && (row * 640 + col) <= 33138) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33139 && (row * 640 + col) <= 33181) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33182 && (row * 640 + col) <= 33194) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33195 && (row * 640 + col) <= 33235) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33236 && (row * 640 + col) <= 33243) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 33244 && (row * 640 + col) <= 33254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33255 && (row * 640 + col) <= 33260) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 33261 && (row * 640 + col) <= 33646) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33647 && (row * 640 + col) <= 33654) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33655 && (row * 640 + col) <= 33680) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33681 && (row * 640 + col) <= 33688) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33689 && (row * 640 + col) <= 33758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33759 && (row * 640 + col) <= 33775) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33776 && (row * 640 + col) <= 33823) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33824 && (row * 640 + col) <= 33835) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33836 && (row * 640 + col) <= 33876) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33877 && (row * 640 + col) <= 33884) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 33885 && (row * 640 + col) <= 33894) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33895 && (row * 640 + col) <= 33900) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 33901 && (row * 640 + col) <= 34286) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34287 && (row * 640 + col) <= 34294) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 34295 && (row * 640 + col) <= 34320) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34321 && (row * 640 + col) <= 34328) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 34329 && (row * 640 + col) <= 34397) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34398 && (row * 640 + col) <= 34413) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 34414 && (row * 640 + col) <= 34464) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34465 && (row * 640 + col) <= 34475) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 34476 && (row * 640 + col) <= 34517) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34518 && (row * 640 + col) <= 34525) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 34526 && (row * 640 + col) <= 34535) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34536 && (row * 640 + col) <= 34541) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 34542 && (row * 640 + col) <= 34927) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34928 && (row * 640 + col) <= 34935) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 34936 && (row * 640 + col) <= 34959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34960 && (row * 640 + col) <= 34968) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 34969 && (row * 640 + col) <= 35036) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35037 && (row * 640 + col) <= 35051) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35052 && (row * 640 + col) <= 35105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35106 && (row * 640 + col) <= 35116) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35117 && (row * 640 + col) <= 35158) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35159 && (row * 640 + col) <= 35166) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 35167 && (row * 640 + col) <= 35175) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35176 && (row * 640 + col) <= 35181) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 35182 && (row * 640 + col) <= 35567) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35568 && (row * 640 + col) <= 35576) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35577 && (row * 640 + col) <= 35599) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35600 && (row * 640 + col) <= 35608) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35609 && (row * 640 + col) <= 35675) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35676 && (row * 640 + col) <= 35689) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35690 && (row * 640 + col) <= 35746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35747 && (row * 640 + col) <= 35756) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35757 && (row * 640 + col) <= 35799) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35800 && (row * 640 + col) <= 35807) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 35808 && (row * 640 + col) <= 35816) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35817 && (row * 640 + col) <= 35821) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 35822 && (row * 640 + col) <= 36207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36208 && (row * 640 + col) <= 36216) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36217 && (row * 640 + col) <= 36238) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36239 && (row * 640 + col) <= 36247) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36248 && (row * 640 + col) <= 36314) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36315 && (row * 640 + col) <= 36327) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36328 && (row * 640 + col) <= 36387) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36388 && (row * 640 + col) <= 36397) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36398 && (row * 640 + col) <= 36440) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36441 && (row * 640 + col) <= 36448) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 36449 && (row * 640 + col) <= 36456) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36457 && (row * 640 + col) <= 36462) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 36463 && (row * 640 + col) <= 36848) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36849 && (row * 640 + col) <= 36857) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36858 && (row * 640 + col) <= 36877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36878 && (row * 640 + col) <= 36887) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36888 && (row * 640 + col) <= 36953) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36954 && (row * 640 + col) <= 36966) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36967 && (row * 640 + col) <= 37028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37029 && (row * 640 + col) <= 37037) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37038 && (row * 640 + col) <= 37081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37082 && (row * 640 + col) <= 37089) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 37090 && (row * 640 + col) <= 37097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37098 && (row * 640 + col) <= 37102) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 37103 && (row * 640 + col) <= 37200) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37201 && (row * 640 + col) <= 37206) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37207 && (row * 640 + col) <= 37488) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37489 && (row * 640 + col) <= 37498) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37499 && (row * 640 + col) <= 37517) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37518 && (row * 640 + col) <= 37526) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37527 && (row * 640 + col) <= 37592) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37593 && (row * 640 + col) <= 37605) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37606 && (row * 640 + col) <= 37668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37669 && (row * 640 + col) <= 37677) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37678 && (row * 640 + col) <= 37722) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37723 && (row * 640 + col) <= 37730) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 37731 && (row * 640 + col) <= 37737) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37738 && (row * 640 + col) <= 37743) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 37744 && (row * 640 + col) <= 37837) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 37838 && (row * 640 + col) <= 37849) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37850 && (row * 640 + col) <= 38129) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38130 && (row * 640 + col) <= 38139) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38140 && (row * 640 + col) <= 38155) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38156 && (row * 640 + col) <= 38166) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38167 && (row * 640 + col) <= 38232) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38233 && (row * 640 + col) <= 38243) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38244 && (row * 640 + col) <= 38309) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38310 && (row * 640 + col) <= 38318) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38319 && (row * 640 + col) <= 38363) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38364 && (row * 640 + col) <= 38370) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 38371 && (row * 640 + col) <= 38377) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38378 && (row * 640 + col) <= 38383) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 38384 && (row * 640 + col) <= 38475) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38476 && (row * 640 + col) <= 38492) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38493 && (row * 640 + col) <= 38769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38770 && (row * 640 + col) <= 38780) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38781 && (row * 640 + col) <= 38794) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38795 && (row * 640 + col) <= 38805) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38806 && (row * 640 + col) <= 38871) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38872 && (row * 640 + col) <= 38882) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38883 && (row * 640 + col) <= 38949) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 38950 && (row * 640 + col) <= 38958) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38959 && (row * 640 + col) <= 39004) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39005 && (row * 640 + col) <= 39011) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 39012 && (row * 640 + col) <= 39017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39018 && (row * 640 + col) <= 39023) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 39024 && (row * 640 + col) <= 39113) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39114 && (row * 640 + col) <= 39134) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39135 && (row * 640 + col) <= 39410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39411 && (row * 640 + col) <= 39422) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39423 && (row * 640 + col) <= 39432) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39433 && (row * 640 + col) <= 39445) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39446 && (row * 640 + col) <= 39510) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39511 && (row * 640 + col) <= 39521) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39522 && (row * 640 + col) <= 39589) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39590 && (row * 640 + col) <= 39598) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39599 && (row * 640 + col) <= 39645) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39646 && (row * 640 + col) <= 39652) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 39653 && (row * 640 + col) <= 39658) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39659 && (row * 640 + col) <= 39663) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 39664 && (row * 640 + col) <= 39750) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 39751 && (row * 640 + col) <= 39777) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39778 && (row * 640 + col) <= 40051) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40052 && (row * 640 + col) <= 40084) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40085 && (row * 640 + col) <= 40150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40151 && (row * 640 + col) <= 40160) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40161 && (row * 640 + col) <= 40229) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40230 && (row * 640 + col) <= 40238) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40239 && (row * 640 + col) <= 40286) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40287 && (row * 640 + col) <= 40293) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 40294 && (row * 640 + col) <= 40298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40299 && (row * 640 + col) <= 40304) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 40305 && (row * 640 + col) <= 40388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40389 && (row * 640 + col) <= 40419) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40420 && (row * 640 + col) <= 40692) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40693 && (row * 640 + col) <= 40723) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40724 && (row * 640 + col) <= 40789) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40790 && (row * 640 + col) <= 40799) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40800 && (row * 640 + col) <= 40869) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40870 && (row * 640 + col) <= 40878) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40879 && (row * 640 + col) <= 40927) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40928 && (row * 640 + col) <= 40934) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 40935 && (row * 640 + col) <= 40938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 40939 && (row * 640 + col) <= 40944) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 40945 && (row * 640 + col) <= 41025) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41026 && (row * 640 + col) <= 41061) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 41062 && (row * 640 + col) <= 41333) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41334 && (row * 640 + col) <= 41362) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 41363 && (row * 640 + col) <= 41429) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41430 && (row * 640 + col) <= 41439) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 41440 && (row * 640 + col) <= 41509) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41510 && (row * 640 + col) <= 41518) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 41519 && (row * 640 + col) <= 41568) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41569 && (row * 640 + col) <= 41575) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 41576 && (row * 640 + col) <= 41578) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41579 && (row * 640 + col) <= 41584) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 41585 && (row * 640 + col) <= 41663) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41664 && (row * 640 + col) <= 41704) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 41705 && (row * 640 + col) <= 41974) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 41975 && (row * 640 + col) <= 42001) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42002 && (row * 640 + col) <= 42069) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42070 && (row * 640 + col) <= 42078) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42079 && (row * 640 + col) <= 42149) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42150 && (row * 640 + col) <= 42158) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42159 && (row * 640 + col) <= 42208) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42209 && (row * 640 + col) <= 42223) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 42224 && (row * 640 + col) <= 42301) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42302 && (row * 640 + col) <= 42346) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42347 && (row * 640 + col) <= 42615) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42616 && (row * 640 + col) <= 42640) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42641 && (row * 640 + col) <= 42708) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42709 && (row * 640 + col) <= 42717) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42718 && (row * 640 + col) <= 42788) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42789 && (row * 640 + col) <= 42797) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42798 && (row * 640 + col) <= 42849) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42850 && (row * 640 + col) <= 42863) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 42864 && (row * 640 + col) <= 42938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 42939 && (row * 640 + col) <= 42989) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42990 && (row * 640 + col) <= 43119) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43120 && (row * 640 + col) <= 43123) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 43124 && (row * 640 + col) <= 43257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43258 && (row * 640 + col) <= 43278) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43279 && (row * 640 + col) <= 43348) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43349 && (row * 640 + col) <= 43357) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43358 && (row * 640 + col) <= 43428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43429 && (row * 640 + col) <= 43437) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43438 && (row * 640 + col) <= 43490) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43491 && (row * 640 + col) <= 43502) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 43503 && (row * 640 + col) <= 43576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43577 && (row * 640 + col) <= 43602) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43603 && (row * 640 + col) <= 43604) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43605 && (row * 640 + col) <= 43631) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43632 && (row * 640 + col) <= 43756) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43757 && (row * 640 + col) <= 43767) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 43768 && (row * 640 + col) <= 43899) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43900 && (row * 640 + col) <= 43916) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43917 && (row * 640 + col) <= 43988) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 43989 && (row * 640 + col) <= 43997) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43998 && (row * 640 + col) <= 44067) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44068 && (row * 640 + col) <= 44077) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44078 && (row * 640 + col) <= 44131) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44132 && (row * 640 + col) <= 44142) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 44143 && (row * 640 + col) <= 44214) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44215 && (row * 640 + col) <= 44240) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44241 && (row * 640 + col) <= 44247) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44248 && (row * 640 + col) <= 44273) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44274 && (row * 640 + col) <= 44393) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44394 && (row * 640 + col) <= 44409) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 44410 && (row * 640 + col) <= 44541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44542 && (row * 640 + col) <= 44554) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44555 && (row * 640 + col) <= 44627) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44628 && (row * 640 + col) <= 44636) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44637 && (row * 640 + col) <= 44706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44707 && (row * 640 + col) <= 44716) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44717 && (row * 640 + col) <= 44772) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44773 && (row * 640 + col) <= 44780) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 44781 && (row * 640 + col) <= 44851) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44852 && (row * 640 + col) <= 44877) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44878 && (row * 640 + col) <= 44890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 44891 && (row * 640 + col) <= 44916) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 44917 && (row * 640 + col) <= 45031) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45032 && (row * 640 + col) <= 45052) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 45053 && (row * 640 + col) <= 45267) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45268 && (row * 640 + col) <= 45276) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 45277 && (row * 640 + col) <= 45345) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45346 && (row * 640 + col) <= 45356) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 45357 && (row * 640 + col) <= 45414) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45415 && (row * 640 + col) <= 45418) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 45419 && (row * 640 + col) <= 45489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45490 && (row * 640 + col) <= 45515) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 45516 && (row * 640 + col) <= 45532) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45533 && (row * 640 + col) <= 45558) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 45559 && (row * 640 + col) <= 45669) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45670 && (row * 640 + col) <= 45694) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 45695 && (row * 640 + col) <= 45907) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45908 && (row * 640 + col) <= 45916) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 45917 && (row * 640 + col) <= 45983) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 45984 && (row * 640 + col) <= 45996) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 45997 && (row * 640 + col) <= 46126) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46127 && (row * 640 + col) <= 46152) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46153 && (row * 640 + col) <= 46174) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46175 && (row * 640 + col) <= 46200) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46201 && (row * 640 + col) <= 46306) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46307 && (row * 640 + col) <= 46336) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 46337 && (row * 640 + col) <= 46547) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46548 && (row * 640 + col) <= 46556) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46557 && (row * 640 + col) <= 46619) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46620 && (row * 640 + col) <= 46635) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46636 && (row * 640 + col) <= 46764) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46765 && (row * 640 + col) <= 46790) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46791 && (row * 640 + col) <= 46817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46818 && (row * 640 + col) <= 46843) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46844 && (row * 640 + col) <= 46944) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 46945 && (row * 640 + col) <= 46979) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 46980 && (row * 640 + col) <= 47187) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 47188 && (row * 640 + col) <= 47196) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 47197 && (row * 640 + col) <= 47239) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 47240 && (row * 640 + col) <= 47274) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 47275 && (row * 640 + col) <= 47402) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 47403 && (row * 640 + col) <= 47428) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 47429 && (row * 640 + col) <= 47459) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 47460 && (row * 640 + col) <= 47485) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 47486 && (row * 640 + col) <= 47581) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 47582 && (row * 640 + col) <= 47621) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 47622 && (row * 640 + col) <= 47827) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 47828 && (row * 640 + col) <= 47836) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 47837 && (row * 640 + col) <= 47873) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 47874 && (row * 640 + col) <= 47913) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 47914 && (row * 640 + col) <= 48039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48040 && (row * 640 + col) <= 48065) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48066 && (row * 640 + col) <= 48102) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48103 && (row * 640 + col) <= 48128) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48129 && (row * 640 + col) <= 48219) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48220 && (row * 640 + col) <= 48264) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 48265 && (row * 640 + col) <= 48467) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48468 && (row * 640 + col) <= 48476) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48477 && (row * 640 + col) <= 48508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48509 && (row * 640 + col) <= 48553) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48554 && (row * 640 + col) <= 48677) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48678 && (row * 640 + col) <= 48703) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48704 && (row * 640 + col) <= 48744) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48745 && (row * 640 + col) <= 48769) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48770 && (row * 640 + col) <= 48856) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48857 && (row * 640 + col) <= 48879) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 48880 && (row * 640 + col) <= 48884) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 48885 && (row * 640 + col) <= 48906) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 48907 && (row * 640 + col) <= 49107) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49108 && (row * 640 + col) <= 49116) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49117 && (row * 640 + col) <= 49145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49146 && (row * 640 + col) <= 49191) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49192 && (row * 640 + col) <= 49316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49317 && (row * 640 + col) <= 49340) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49341 && (row * 640 + col) <= 49386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49387 && (row * 640 + col) <= 49411) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49412 && (row * 640 + col) <= 49494) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49495 && (row * 640 + col) <= 49517) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 49518 && (row * 640 + col) <= 49526) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49527 && (row * 640 + col) <= 49548) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 49549 && (row * 640 + col) <= 49747) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49748 && (row * 640 + col) <= 49756) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49757 && (row * 640 + col) <= 49782) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49783 && (row * 640 + col) <= 49830) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49831 && (row * 640 + col) <= 49955) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 49956 && (row * 640 + col) <= 49978) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49979 && (row * 640 + col) <= 50029) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50030 && (row * 640 + col) <= 50052) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 50053 && (row * 640 + col) <= 50131) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50132 && (row * 640 + col) <= 50154) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 50155 && (row * 640 + col) <= 50169) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50170 && (row * 640 + col) <= 50191) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 50192 && (row * 640 + col) <= 50388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50389 && (row * 640 + col) <= 50397) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 50398 && (row * 640 + col) <= 50419) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50420 && (row * 640 + col) <= 50468) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 50469 && (row * 640 + col) <= 50594) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50595 && (row * 640 + col) <= 50615) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 50616 && (row * 640 + col) <= 50671) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50672 && (row * 640 + col) <= 50693) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 50694 && (row * 640 + col) <= 50769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50770 && (row * 640 + col) <= 50792) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 50793 && (row * 640 + col) <= 50811) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 50812 && (row * 640 + col) <= 50833) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 50834 && (row * 640 + col) <= 51028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51029 && (row * 640 + col) <= 51037) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51038 && (row * 640 + col) <= 51058) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51059 && (row * 640 + col) <= 51106) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51107 && (row * 640 + col) <= 51233) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51234 && (row * 640 + col) <= 51253) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51254 && (row * 640 + col) <= 51313) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51314 && (row * 640 + col) <= 51334) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51335 && (row * 640 + col) <= 51407) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51408 && (row * 640 + col) <= 51429) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 51430 && (row * 640 + col) <= 51453) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51454 && (row * 640 + col) <= 51475) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 51476 && (row * 640 + col) <= 51668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51669 && (row * 640 + col) <= 51678) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51679 && (row * 640 + col) <= 51695) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51696 && (row * 640 + col) <= 51744) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51745 && (row * 640 + col) <= 51872) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51873 && (row * 640 + col) <= 51890) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51891 && (row * 640 + col) <= 51956) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 51957 && (row * 640 + col) <= 51974) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51975 && (row * 640 + col) <= 52044) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52045 && (row * 640 + col) <= 52067) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 52068 && (row * 640 + col) <= 52096) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52097 && (row * 640 + col) <= 52118) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 52119 && (row * 640 + col) <= 52309) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52310 && (row * 640 + col) <= 52319) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 52320 && (row * 640 + col) <= 52333) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52334 && (row * 640 + col) <= 52369) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 52370 && (row * 640 + col) <= 52511) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52512 && (row * 640 + col) <= 52528) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 52529 && (row * 640 + col) <= 52598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52599 && (row * 640 + col) <= 52615) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 52616 && (row * 640 + col) <= 52682) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52683 && (row * 640 + col) <= 52705) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 52706 && (row * 640 + col) <= 52738) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52739 && (row * 640 + col) <= 52760) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 52761 && (row * 640 + col) <= 52949) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52950 && (row * 640 + col) <= 52960) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 52961 && (row * 640 + col) <= 52971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 52972 && (row * 640 + col) <= 52997) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 52998 && (row * 640 + col) <= 53151) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53152 && (row * 640 + col) <= 53165) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53166 && (row * 640 + col) <= 53241) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53242 && (row * 640 + col) <= 53256) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53257 && (row * 640 + col) <= 53320) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53321 && (row * 640 + col) <= 53342) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 53343 && (row * 640 + col) <= 53381) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53382 && (row * 640 + col) <= 53402) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 53403 && (row * 640 + col) <= 53590) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53591 && (row * 640 + col) <= 53604) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53605 && (row * 640 + col) <= 53606) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53607 && (row * 640 + col) <= 53631) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53632 && (row * 640 + col) <= 53791) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53792 && (row * 640 + col) <= 53803) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53804 && (row * 640 + col) <= 53883) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53884 && (row * 640 + col) <= 53896) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53897 && (row * 640 + col) <= 53959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 53960 && (row * 640 + col) <= 53980) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 53981 && (row * 640 + col) <= 54023) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54024 && (row * 640 + col) <= 54043) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 54044 && (row * 640 + col) <= 54230) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54231 && (row * 640 + col) <= 54268) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 54269 && (row * 640 + col) <= 54430) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54431 && (row * 640 + col) <= 54442) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 54443 && (row * 640 + col) <= 54525) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54526 && (row * 640 + col) <= 54537) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 54538 && (row * 640 + col) <= 54598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54599 && (row * 640 + col) <= 54618) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 54619 && (row * 640 + col) <= 54665) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54666 && (row * 640 + col) <= 54684) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 54685 && (row * 640 + col) <= 54871) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54872 && (row * 640 + col) <= 54905) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 54906 && (row * 640 + col) <= 54992) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 54993 && (row * 640 + col) <= 55003) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55004 && (row * 640 + col) <= 55070) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55071 && (row * 640 + col) <= 55081) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55082 && (row * 640 + col) <= 55166) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55167 && (row * 640 + col) <= 55177) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55178 && (row * 640 + col) <= 55237) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55238 && (row * 640 + col) <= 55255) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 55256 && (row * 640 + col) <= 55308) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55309 && (row * 640 + col) <= 55325) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 55326 && (row * 640 + col) <= 55512) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55513 && (row * 640 + col) <= 55543) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55544 && (row * 640 + col) <= 55629) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55630 && (row * 640 + col) <= 55646) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55647 && (row * 640 + col) <= 55709) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55710 && (row * 640 + col) <= 55720) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55721 && (row * 640 + col) <= 55806) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55807 && (row * 640 + col) <= 55817) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55818 && (row * 640 + col) <= 55876) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55877 && (row * 640 + col) <= 55893) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 55894 && (row * 640 + col) <= 55950) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 55951 && (row * 640 + col) <= 55966) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 55967 && (row * 640 + col) <= 56153) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56154 && (row * 640 + col) <= 56181) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 56182 && (row * 640 + col) <= 56267) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56268 && (row * 640 + col) <= 56288) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 56289 && (row * 640 + col) <= 56349) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56350 && (row * 640 + col) <= 56360) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 56361 && (row * 640 + col) <= 56447) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56448 && (row * 640 + col) <= 56458) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 56459 && (row * 640 + col) <= 56516) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56517 && (row * 640 + col) <= 56530) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 56531 && (row * 640 + col) <= 56593) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56594 && (row * 640 + col) <= 56607) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 56608 && (row * 640 + col) <= 56794) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56795 && (row * 640 + col) <= 56819) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 56820 && (row * 640 + col) <= 56906) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56907 && (row * 640 + col) <= 56930) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 56931 && (row * 640 + col) <= 56989) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56990 && (row * 640 + col) <= 56999) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57000 && (row * 640 + col) <= 57087) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57088 && (row * 640 + col) <= 57098) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57099 && (row * 640 + col) <= 57155) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57156 && (row * 640 + col) <= 57168) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 57169 && (row * 640 + col) <= 57235) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57236 && (row * 640 + col) <= 57247) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 57248 && (row * 640 + col) <= 57435) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57436 && (row * 640 + col) <= 57456) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57457 && (row * 640 + col) <= 57544) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57545 && (row * 640 + col) <= 57572) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57573 && (row * 640 + col) <= 57628) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57629 && (row * 640 + col) <= 57639) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57640 && (row * 640 + col) <= 57728) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57729 && (row * 640 + col) <= 57739) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57740 && (row * 640 + col) <= 57795) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57796 && (row * 640 + col) <= 57806) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 57807 && (row * 640 + col) <= 57877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57878 && (row * 640 + col) <= 57887) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 57888 && (row * 640 + col) <= 58077) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58078 && (row * 640 + col) <= 58094) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58095 && (row * 640 + col) <= 58184) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58185 && (row * 640 + col) <= 58213) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58214 && (row * 640 + col) <= 58268) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58269 && (row * 640 + col) <= 58278) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58279 && (row * 640 + col) <= 58368) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58369 && (row * 640 + col) <= 58379) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58380 && (row * 640 + col) <= 58435) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58436 && (row * 640 + col) <= 58444) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 58445 && (row * 640 + col) <= 58518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58519 && (row * 640 + col) <= 58528) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 58529 && (row * 640 + col) <= 58720) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58721 && (row * 640 + col) <= 58730) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58731 && (row * 640 + col) <= 58823) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58824 && (row * 640 + col) <= 58854) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58855 && (row * 640 + col) <= 58907) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58908 && (row * 640 + col) <= 58918) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58919 && (row * 640 + col) <= 59009) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59010 && (row * 640 + col) <= 59019) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 59020 && (row * 640 + col) <= 59074) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59075 && (row * 640 + col) <= 59084) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 59085 && (row * 640 + col) <= 59159) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59160 && (row * 640 + col) <= 59168) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 59169 && (row * 640 + col) <= 59462) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59463 && (row * 640 + col) <= 59495) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 59496 && (row * 640 + col) <= 59547) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59548 && (row * 640 + col) <= 59558) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 59559 && (row * 640 + col) <= 59649) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59650 && (row * 640 + col) <= 59660) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 59661 && (row * 640 + col) <= 59714) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59715 && (row * 640 + col) <= 59723) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 59724 && (row * 640 + col) <= 59799) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59800 && (row * 640 + col) <= 59809) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 59810 && (row * 640 + col) <= 60101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60102 && (row * 640 + col) <= 60116) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60117 && (row * 640 + col) <= 60119) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60120 && (row * 640 + col) <= 60136) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60137 && (row * 640 + col) <= 60186) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60187 && (row * 640 + col) <= 60197) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60198 && (row * 640 + col) <= 60289) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60290 && (row * 640 + col) <= 60300) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60301 && (row * 640 + col) <= 60353) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60354 && (row * 640 + col) <= 60363) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 60364 && (row * 640 + col) <= 60440) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60441 && (row * 640 + col) <= 60449) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 60450 && (row * 640 + col) <= 60741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60742 && (row * 640 + col) <= 60752) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60753 && (row * 640 + col) <= 60763) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60764 && (row * 640 + col) <= 60777) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60778 && (row * 640 + col) <= 60826) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60827 && (row * 640 + col) <= 60837) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60838 && (row * 640 + col) <= 60930) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60931 && (row * 640 + col) <= 60941) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60942 && (row * 640 + col) <= 60993) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60994 && (row * 640 + col) <= 61002) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 61003 && (row * 640 + col) <= 61080) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61081 && (row * 640 + col) <= 61090) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 61091 && (row * 640 + col) <= 61380) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61381 && (row * 640 + col) <= 61391) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 61392 && (row * 640 + col) <= 61405) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61406 && (row * 640 + col) <= 61418) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 61419 && (row * 640 + col) <= 61466) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61467 && (row * 640 + col) <= 61476) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 61477 && (row * 640 + col) <= 61570) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61571 && (row * 640 + col) <= 61581) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 61582 && (row * 640 + col) <= 61632) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61633 && (row * 640 + col) <= 61642) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 61643 && (row * 640 + col) <= 61721) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61722 && (row * 640 + col) <= 61730) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 61731 && (row * 640 + col) <= 62020) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62021 && (row * 640 + col) <= 62030) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62031 && (row * 640 + col) <= 62047) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62048 && (row * 640 + col) <= 62059) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62060 && (row * 640 + col) <= 62105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62106 && (row * 640 + col) <= 62116) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62117 && (row * 640 + col) <= 62211) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62212 && (row * 640 + col) <= 62222) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62223 && (row * 640 + col) <= 62272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62273 && (row * 640 + col) <= 62282) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 62283 && (row * 640 + col) <= 62361) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62362 && (row * 640 + col) <= 62370) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 62371 && (row * 640 + col) <= 62598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62599 && (row * 640 + col) <= 62614) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 62615 && (row * 640 + col) <= 62659) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62660 && (row * 640 + col) <= 62669) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62670 && (row * 640 + col) <= 62688) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62689 && (row * 640 + col) <= 62699) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62700 && (row * 640 + col) <= 62745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62746 && (row * 640 + col) <= 62756) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62757 && (row * 640 + col) <= 62851) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62852 && (row * 640 + col) <= 62862) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62863 && (row * 640 + col) <= 62912) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62913 && (row * 640 + col) <= 62921) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 62922 && (row * 640 + col) <= 63002) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63003 && (row * 640 + col) <= 63011) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 63012 && (row * 640 + col) <= 63234) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63235 && (row * 640 + col) <= 63258) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 63259 && (row * 640 + col) <= 63299) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63300 && (row * 640 + col) <= 63308) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63309 && (row * 640 + col) <= 63329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63330 && (row * 640 + col) <= 63340) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63341 && (row * 640 + col) <= 63384) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63385 && (row * 640 + col) <= 63395) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63396 && (row * 640 + col) <= 63491) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63492 && (row * 640 + col) <= 63502) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63503 && (row * 640 + col) <= 63551) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63552 && (row * 640 + col) <= 63561) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 63562 && (row * 640 + col) <= 63642) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63643 && (row * 640 + col) <= 63651) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 63652 && (row * 640 + col) <= 63714) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63715 && (row * 640 + col) <= 63731) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63732 && (row * 640 + col) <= 63871) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63872 && (row * 640 + col) <= 63901) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 63902 && (row * 640 + col) <= 63939) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63940 && (row * 640 + col) <= 63948) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63949 && (row * 640 + col) <= 63970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63971 && (row * 640 + col) <= 63981) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63982 && (row * 640 + col) <= 64024) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64025 && (row * 640 + col) <= 64035) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64036 && (row * 640 + col) <= 64132) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64133 && (row * 640 + col) <= 64143) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64144 && (row * 640 + col) <= 64191) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64192 && (row * 640 + col) <= 64200) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 64201 && (row * 640 + col) <= 64282) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64283 && (row * 640 + col) <= 64292) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 64293 && (row * 640 + col) <= 64353) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64354 && (row * 640 + col) <= 64373) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64374 && (row * 640 + col) <= 64509) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64510 && (row * 640 + col) <= 64543) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 64544 && (row * 640 + col) <= 64579) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64580 && (row * 640 + col) <= 64588) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64589 && (row * 640 + col) <= 64611) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64612 && (row * 640 + col) <= 64621) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64622 && (row * 640 + col) <= 64664) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64665 && (row * 640 + col) <= 64674) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64675 && (row * 640 + col) <= 64772) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64773 && (row * 640 + col) <= 64783) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64784 && (row * 640 + col) <= 64830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64831 && (row * 640 + col) <= 64840) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 64841 && (row * 640 + col) <= 64923) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64924 && (row * 640 + col) <= 64932) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 64933 && (row * 640 + col) <= 64992) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64993 && (row * 640 + col) <= 65014) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65015 && (row * 640 + col) <= 65147) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65148 && (row * 640 + col) <= 65185) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 65186 && (row * 640 + col) <= 65219) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65220 && (row * 640 + col) <= 65227) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65228 && (row * 640 + col) <= 65252) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65253 && (row * 640 + col) <= 65262) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65263 && (row * 640 + col) <= 65303) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65304 && (row * 640 + col) <= 65314) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65315 && (row * 640 + col) <= 65413) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65414 && (row * 640 + col) <= 65424) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65425 && (row * 640 + col) <= 65470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65471 && (row * 640 + col) <= 65480) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 65481 && (row * 640 + col) <= 65563) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65564 && (row * 640 + col) <= 65572) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 65573 && (row * 640 + col) <= 65631) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65632 && (row * 640 + col) <= 65655) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65656 && (row * 640 + col) <= 65785) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65786 && (row * 640 + col) <= 65827) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 65828 && (row * 640 + col) <= 65859) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65860 && (row * 640 + col) <= 65867) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65868 && (row * 640 + col) <= 65892) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65893 && (row * 640 + col) <= 65902) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65903 && (row * 640 + col) <= 65943) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65944 && (row * 640 + col) <= 65954) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65955 && (row * 640 + col) <= 66053) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66054 && (row * 640 + col) <= 66064) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66065 && (row * 640 + col) <= 66110) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66111 && (row * 640 + col) <= 66119) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 66120 && (row * 640 + col) <= 66204) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66205 && (row * 640 + col) <= 66213) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 66214 && (row * 640 + col) <= 66270) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66271 && (row * 640 + col) <= 66295) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66296 && (row * 640 + col) <= 66423) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66424 && (row * 640 + col) <= 66469) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 66470 && (row * 640 + col) <= 66499) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66500 && (row * 640 + col) <= 66507) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66508 && (row * 640 + col) <= 66533) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66534 && (row * 640 + col) <= 66543) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66544 && (row * 640 + col) <= 66582) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66583 && (row * 640 + col) <= 66593) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66594 && (row * 640 + col) <= 66694) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66695 && (row * 640 + col) <= 66704) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66705 && (row * 640 + col) <= 66749) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66750 && (row * 640 + col) <= 66759) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 66760 && (row * 640 + col) <= 66844) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66845 && (row * 640 + col) <= 66853) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 66854 && (row * 640 + col) <= 66910) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66911 && (row * 640 + col) <= 66917) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66918 && (row * 640 + col) <= 66929) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66930 && (row * 640 + col) <= 66936) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66937 && (row * 640 + col) <= 67062) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67063 && (row * 640 + col) <= 67110) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 67111 && (row * 640 + col) <= 67139) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67140 && (row * 640 + col) <= 67147) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67148 && (row * 640 + col) <= 67174) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67175 && (row * 640 + col) <= 67183) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67184 && (row * 640 + col) <= 67222) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67223 && (row * 640 + col) <= 67233) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67234 && (row * 640 + col) <= 67334) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67335 && (row * 640 + col) <= 67345) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67346 && (row * 640 + col) <= 67389) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67390 && (row * 640 + col) <= 67398) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 67399 && (row * 640 + col) <= 67484) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67485 && (row * 640 + col) <= 67494) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 67495 && (row * 640 + col) <= 67549) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67550 && (row * 640 + col) <= 67555) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67556 && (row * 640 + col) <= 67570) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67571 && (row * 640 + col) <= 67576) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67577 && (row * 640 + col) <= 67700) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67701 && (row * 640 + col) <= 67752) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 67753 && (row * 640 + col) <= 67779) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67780 && (row * 640 + col) <= 67788) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67789 && (row * 640 + col) <= 67814) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67815 && (row * 640 + col) <= 67824) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67825 && (row * 640 + col) <= 67861) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67862 && (row * 640 + col) <= 67872) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67873 && (row * 640 + col) <= 67974) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67975 && (row * 640 + col) <= 67985) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67986 && (row * 640 + col) <= 68028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68029 && (row * 640 + col) <= 68038) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 68039 && (row * 640 + col) <= 68125) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68126 && (row * 640 + col) <= 68134) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 68135 && (row * 640 + col) <= 68189) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68190 && (row * 640 + col) <= 68195) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68196 && (row * 640 + col) <= 68211) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68212 && (row * 640 + col) <= 68217) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68218 && (row * 640 + col) <= 68339) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68340 && (row * 640 + col) <= 68362) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 68363 && (row * 640 + col) <= 68370) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68371 && (row * 640 + col) <= 68393) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 68394 && (row * 640 + col) <= 68419) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68420 && (row * 640 + col) <= 68428) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68429 && (row * 640 + col) <= 68455) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68456 && (row * 640 + col) <= 68464) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68465 && (row * 640 + col) <= 68501) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68502 && (row * 640 + col) <= 68512) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68513 && (row * 640 + col) <= 68615) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68616 && (row * 640 + col) <= 68625) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68626 && (row * 640 + col) <= 68668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68669 && (row * 640 + col) <= 68677) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 68678 && (row * 640 + col) <= 68765) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68766 && (row * 640 + col) <= 68775) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 68776 && (row * 640 + col) <= 68829) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68830 && (row * 640 + col) <= 68834) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68835 && (row * 640 + col) <= 68851) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68852 && (row * 640 + col) <= 68857) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68858 && (row * 640 + col) <= 68978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68979 && (row * 640 + col) <= 68996) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 68997 && (row * 640 + col) <= 69016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69017 && (row * 640 + col) <= 69034) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 69035 && (row * 640 + col) <= 69059) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69060 && (row * 640 + col) <= 69068) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69069 && (row * 640 + col) <= 69095) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69096 && (row * 640 + col) <= 69105) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69106 && (row * 640 + col) <= 69141) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69142 && (row * 640 + col) <= 69151) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69152 && (row * 640 + col) <= 69255) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69256 && (row * 640 + col) <= 69266) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69267 && (row * 640 + col) <= 69307) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69308 && (row * 640 + col) <= 69317) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 69318 && (row * 640 + col) <= 69406) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69407 && (row * 640 + col) <= 69415) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 69416 && (row * 640 + col) <= 69469) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69470 && (row * 640 + col) <= 69474) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69475 && (row * 640 + col) <= 69491) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69492 && (row * 640 + col) <= 69497) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69498 && (row * 640 + col) <= 69617) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69618 && (row * 640 + col) <= 69634) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 69635 && (row * 640 + col) <= 69658) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69659 && (row * 640 + col) <= 69675) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 69676 && (row * 640 + col) <= 69699) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69700 && (row * 640 + col) <= 69708) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69709 && (row * 640 + col) <= 69736) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69737 && (row * 640 + col) <= 69745) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69746 && (row * 640 + col) <= 69780) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69781 && (row * 640 + col) <= 69791) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69792 && (row * 640 + col) <= 69896) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69897 && (row * 640 + col) <= 69906) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69907 && (row * 640 + col) <= 69947) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69948 && (row * 640 + col) <= 69957) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 69958 && (row * 640 + col) <= 70046) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70047 && (row * 640 + col) <= 70055) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 70056 && (row * 640 + col) <= 70109) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70110 && (row * 640 + col) <= 70114) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70115 && (row * 640 + col) <= 70131) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70132 && (row * 640 + col) <= 70137) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70138 && (row * 640 + col) <= 70256) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70257 && (row * 640 + col) <= 70272) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 70273 && (row * 640 + col) <= 70300) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70301 && (row * 640 + col) <= 70316) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 70317 && (row * 640 + col) <= 70340) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70341 && (row * 640 + col) <= 70349) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70350 && (row * 640 + col) <= 70376) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70377 && (row * 640 + col) <= 70385) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70386 && (row * 640 + col) <= 70420) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70421 && (row * 640 + col) <= 70431) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70432 && (row * 640 + col) <= 70536) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70537 && (row * 640 + col) <= 70547) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70548 && (row * 640 + col) <= 70587) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70588 && (row * 640 + col) <= 70596) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 70597 && (row * 640 + col) <= 70687) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70688 && (row * 640 + col) <= 70696) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 70697 && (row * 640 + col) <= 70749) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70750 && (row * 640 + col) <= 70754) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70755 && (row * 640 + col) <= 70771) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70772 && (row * 640 + col) <= 70777) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70778 && (row * 640 + col) <= 70895) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70896 && (row * 640 + col) <= 70910) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 70911 && (row * 640 + col) <= 70942) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70943 && (row * 640 + col) <= 70957) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 70958 && (row * 640 + col) <= 70980) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70981 && (row * 640 + col) <= 70989) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70990 && (row * 640 + col) <= 71017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71018 && (row * 640 + col) <= 71026) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71027 && (row * 640 + col) <= 71059) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71060 && (row * 640 + col) <= 71070) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71071 && (row * 640 + col) <= 71176) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71177 && (row * 640 + col) <= 71187) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71188 && (row * 640 + col) <= 71226) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71227 && (row * 640 + col) <= 71236) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 71237 && (row * 640 + col) <= 71327) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71328 && (row * 640 + col) <= 71336) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 71337 && (row * 640 + col) <= 71389) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71390 && (row * 640 + col) <= 71394) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71395 && (row * 640 + col) <= 71411) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71412 && (row * 640 + col) <= 71417) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71418 && (row * 640 + col) <= 71534) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71535 && (row * 640 + col) <= 71548) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 71549 && (row * 640 + col) <= 71584) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71585 && (row * 640 + col) <= 71598) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 71599 && (row * 640 + col) <= 71620) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71621 && (row * 640 + col) <= 71630) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71631 && (row * 640 + col) <= 71657) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71658 && (row * 640 + col) <= 71666) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71667 && (row * 640 + col) <= 71699) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71700 && (row * 640 + col) <= 71710) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71711 && (row * 640 + col) <= 71817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71818 && (row * 640 + col) <= 71828) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71829 && (row * 640 + col) <= 71866) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71867 && (row * 640 + col) <= 71875) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 71876 && (row * 640 + col) <= 71967) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71968 && (row * 640 + col) <= 71977) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 71978 && (row * 640 + col) <= 72029) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72030 && (row * 640 + col) <= 72034) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72035 && (row * 640 + col) <= 72051) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72052 && (row * 640 + col) <= 72057) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72058 && (row * 640 + col) <= 72173) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72174 && (row * 640 + col) <= 72187) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 72188 && (row * 640 + col) <= 72225) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72226 && (row * 640 + col) <= 72239) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 72240 && (row * 640 + col) <= 72261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72262 && (row * 640 + col) <= 72270) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72271 && (row * 640 + col) <= 72297) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72298 && (row * 640 + col) <= 72307) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72308 && (row * 640 + col) <= 72338) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72339 && (row * 640 + col) <= 72349) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72350 && (row * 640 + col) <= 72457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72458 && (row * 640 + col) <= 72468) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72469 && (row * 640 + col) <= 72505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72506 && (row * 640 + col) <= 72515) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 72516 && (row * 640 + col) <= 72608) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72609 && (row * 640 + col) <= 72617) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 72618 && (row * 640 + col) <= 72669) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72670 && (row * 640 + col) <= 72674) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72675 && (row * 640 + col) <= 72691) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72692 && (row * 640 + col) <= 72697) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72698 && (row * 640 + col) <= 72812) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72813 && (row * 640 + col) <= 72825) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 72826 && (row * 640 + col) <= 72867) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72868 && (row * 640 + col) <= 72880) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 72881 && (row * 640 + col) <= 72901) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72902 && (row * 640 + col) <= 72910) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72911 && (row * 640 + col) <= 72938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72939 && (row * 640 + col) <= 72947) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72948 && (row * 640 + col) <= 72978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72979 && (row * 640 + col) <= 72989) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72990 && (row * 640 + col) <= 73097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73098 && (row * 640 + col) <= 73108) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73109 && (row * 640 + col) <= 73145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73146 && (row * 640 + col) <= 73155) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 73156 && (row * 640 + col) <= 73248) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73249 && (row * 640 + col) <= 73257) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 73258 && (row * 640 + col) <= 73309) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73310 && (row * 640 + col) <= 73314) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73315 && (row * 640 + col) <= 73331) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73332 && (row * 640 + col) <= 73337) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73338 && (row * 640 + col) <= 73452) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73453 && (row * 640 + col) <= 73464) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 73465 && (row * 640 + col) <= 73508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73509 && (row * 640 + col) <= 73520) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 73521 && (row * 640 + col) <= 73541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73542 && (row * 640 + col) <= 73551) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73552 && (row * 640 + col) <= 73578) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73579 && (row * 640 + col) <= 73587) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73588 && (row * 640 + col) <= 73618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73619 && (row * 640 + col) <= 73629) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73630 && (row * 640 + col) <= 73738) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73739 && (row * 640 + col) <= 73749) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73750 && (row * 640 + col) <= 73785) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73786 && (row * 640 + col) <= 73794) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 73795 && (row * 640 + col) <= 73889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73890 && (row * 640 + col) <= 73898) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 73899 && (row * 640 + col) <= 73949) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73950 && (row * 640 + col) <= 73954) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73955 && (row * 640 + col) <= 73971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73972 && (row * 640 + col) <= 73977) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73978 && (row * 640 + col) <= 74091) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74092 && (row * 640 + col) <= 74103) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 74104 && (row * 640 + col) <= 74149) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74150 && (row * 640 + col) <= 74161) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 74162 && (row * 640 + col) <= 74182) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74183 && (row * 640 + col) <= 74191) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74192 && (row * 640 + col) <= 74218) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74219 && (row * 640 + col) <= 74227) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74228 && (row * 640 + col) <= 74257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74258 && (row * 640 + col) <= 74268) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74269 && (row * 640 + col) <= 74378) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74379 && (row * 640 + col) <= 74389) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74390 && (row * 640 + col) <= 74424) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74425 && (row * 640 + col) <= 74434) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 74435 && (row * 640 + col) <= 74529) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74530 && (row * 640 + col) <= 74538) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 74539 && (row * 640 + col) <= 74589) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74590 && (row * 640 + col) <= 74594) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74595 && (row * 640 + col) <= 74611) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74612 && (row * 640 + col) <= 74617) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74618 && (row * 640 + col) <= 74730) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74731 && (row * 640 + col) <= 74742) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 74743 && (row * 640 + col) <= 74790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74791 && (row * 640 + col) <= 74802) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 74803 && (row * 640 + col) <= 74822) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74823 && (row * 640 + col) <= 74832) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74833 && (row * 640 + col) <= 74859) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74860 && (row * 640 + col) <= 74868) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74869 && (row * 640 + col) <= 74897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74898 && (row * 640 + col) <= 74908) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74909 && (row * 640 + col) <= 75019) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75020 && (row * 640 + col) <= 75030) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75031 && (row * 640 + col) <= 75064) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75065 && (row * 640 + col) <= 75073) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 75074 && (row * 640 + col) <= 75169) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75170 && (row * 640 + col) <= 75179) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 75180 && (row * 640 + col) <= 75229) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75230 && (row * 640 + col) <= 75234) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75235 && (row * 640 + col) <= 75251) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75252 && (row * 640 + col) <= 75257) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75258 && (row * 640 + col) <= 75370) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75371 && (row * 640 + col) <= 75381) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 75382 && (row * 640 + col) <= 75431) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75432 && (row * 640 + col) <= 75442) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 75443 && (row * 640 + col) <= 75463) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75464 && (row * 640 + col) <= 75472) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75473 && (row * 640 + col) <= 75499) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75500 && (row * 640 + col) <= 75508) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75509 && (row * 640 + col) <= 75536) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75537 && (row * 640 + col) <= 75547) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75548 && (row * 640 + col) <= 75659) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75660 && (row * 640 + col) <= 75670) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75671 && (row * 640 + col) <= 75703) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75704 && (row * 640 + col) <= 75713) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 75714 && (row * 640 + col) <= 75810) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75811 && (row * 640 + col) <= 75819) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 75820 && (row * 640 + col) <= 75869) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75870 && (row * 640 + col) <= 75874) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75875 && (row * 640 + col) <= 75891) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75892 && (row * 640 + col) <= 75897) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75898 && (row * 640 + col) <= 76009) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76010 && (row * 640 + col) <= 76020) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 76021 && (row * 640 + col) <= 76072) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76073 && (row * 640 + col) <= 76083) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 76084 && (row * 640 + col) <= 76103) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76104 && (row * 640 + col) <= 76113) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76114 && (row * 640 + col) <= 76139) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76140 && (row * 640 + col) <= 76148) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76149 && (row * 640 + col) <= 76176) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76177 && (row * 640 + col) <= 76187) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76188 && (row * 640 + col) <= 76299) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76300 && (row * 640 + col) <= 76310) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76311 && (row * 640 + col) <= 76343) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76344 && (row * 640 + col) <= 76352) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 76353 && (row * 640 + col) <= 76450) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76451 && (row * 640 + col) <= 76459) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 76460 && (row * 640 + col) <= 76509) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76510 && (row * 640 + col) <= 76514) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76515 && (row * 640 + col) <= 76531) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76532 && (row * 640 + col) <= 76537) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76538 && (row * 640 + col) <= 76649) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76650 && (row * 640 + col) <= 76660) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 76661 && (row * 640 + col) <= 76712) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76713 && (row * 640 + col) <= 76723) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 76724 && (row * 640 + col) <= 76744) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76745 && (row * 640 + col) <= 76753) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76754 && (row * 640 + col) <= 76779) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76780 && (row * 640 + col) <= 76788) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76789 && (row * 640 + col) <= 76816) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76817 && (row * 640 + col) <= 76826) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76827 && (row * 640 + col) <= 76940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76941 && (row * 640 + col) <= 76951) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76952 && (row * 640 + col) <= 76982) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76983 && (row * 640 + col) <= 76992) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 76993 && (row * 640 + col) <= 77091) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77092 && (row * 640 + col) <= 77100) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 77101 && (row * 640 + col) <= 77149) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77150 && (row * 640 + col) <= 77154) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77155 && (row * 640 + col) <= 77171) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77172 && (row * 640 + col) <= 77177) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77178 && (row * 640 + col) <= 77288) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77289 && (row * 640 + col) <= 77299) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 77300 && (row * 640 + col) <= 77353) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77354 && (row * 640 + col) <= 77364) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 77365 && (row * 640 + col) <= 77384) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77385 && (row * 640 + col) <= 77393) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77394 && (row * 640 + col) <= 77420) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77421 && (row * 640 + col) <= 77429) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77430 && (row * 640 + col) <= 77455) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77456 && (row * 640 + col) <= 77466) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77467 && (row * 640 + col) <= 77580) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77581 && (row * 640 + col) <= 77591) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77592 && (row * 640 + col) <= 77622) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77623 && (row * 640 + col) <= 77632) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 77633 && (row * 640 + col) <= 77731) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77732 && (row * 640 + col) <= 77740) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 77741 && (row * 640 + col) <= 77789) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77790 && (row * 640 + col) <= 77794) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77795 && (row * 640 + col) <= 77811) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77812 && (row * 640 + col) <= 77816) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77817 && (row * 640 + col) <= 77928) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77929 && (row * 640 + col) <= 77938) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 77939 && (row * 640 + col) <= 77994) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77995 && (row * 640 + col) <= 78004) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 78005 && (row * 640 + col) <= 78024) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78025 && (row * 640 + col) <= 78034) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78035 && (row * 640 + col) <= 78060) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78061 && (row * 640 + col) <= 78069) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78070 && (row * 640 + col) <= 78095) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78096 && (row * 640 + col) <= 78106) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78107 && (row * 640 + col) <= 78221) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78222 && (row * 640 + col) <= 78232) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78233 && (row * 640 + col) <= 78262) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78263 && (row * 640 + col) <= 78271) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 78272 && (row * 640 + col) <= 78372) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78373 && (row * 640 + col) <= 78381) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 78382 && (row * 640 + col) <= 78429) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78430 && (row * 640 + col) <= 78434) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78435 && (row * 640 + col) <= 78451) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78452 && (row * 640 + col) <= 78456) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78457 && (row * 640 + col) <= 78567) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78568 && (row * 640 + col) <= 78578) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 78579 && (row * 640 + col) <= 78634) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78635 && (row * 640 + col) <= 78645) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 78646 && (row * 640 + col) <= 78665) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78666 && (row * 640 + col) <= 78674) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78675 && (row * 640 + col) <= 78700) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78701 && (row * 640 + col) <= 78709) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78710 && (row * 640 + col) <= 78735) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78736 && (row * 640 + col) <= 78745) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78746 && (row * 640 + col) <= 78861) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78862 && (row * 640 + col) <= 78872) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78873 && (row * 640 + col) <= 78901) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78902 && (row * 640 + col) <= 78911) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 78912 && (row * 640 + col) <= 79012) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79013 && (row * 640 + col) <= 79021) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 79022 && (row * 640 + col) <= 79069) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79070 && (row * 640 + col) <= 79075) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79076 && (row * 640 + col) <= 79091) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79092 && (row * 640 + col) <= 79096) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79097 && (row * 640 + col) <= 79207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79208 && (row * 640 + col) <= 79217) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 79218 && (row * 640 + col) <= 79275) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79276 && (row * 640 + col) <= 79285) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 79286 && (row * 640 + col) <= 79305) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79306 && (row * 640 + col) <= 79314) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79315 && (row * 640 + col) <= 79340) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79341 && (row * 640 + col) <= 79349) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79350 && (row * 640 + col) <= 79374) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79375 && (row * 640 + col) <= 79385) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79386 && (row * 640 + col) <= 79502) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79503 && (row * 640 + col) <= 79512) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79513 && (row * 640 + col) <= 79541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79542 && (row * 640 + col) <= 79550) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 79551 && (row * 640 + col) <= 79652) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79653 && (row * 640 + col) <= 79661) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 79662 && (row * 640 + col) <= 79709) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79710 && (row * 640 + col) <= 79716) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79717 && (row * 640 + col) <= 79730) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79731 && (row * 640 + col) <= 79736) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79737 && (row * 640 + col) <= 79847) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79848 && (row * 640 + col) <= 79857) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 79858 && (row * 640 + col) <= 79915) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79916 && (row * 640 + col) <= 79926) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 79927 && (row * 640 + col) <= 79945) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79946 && (row * 640 + col) <= 79955) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79956 && (row * 640 + col) <= 79981) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79982 && (row * 640 + col) <= 79989) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79990 && (row * 640 + col) <= 80014) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80015 && (row * 640 + col) <= 80024) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80025 && (row * 640 + col) <= 80142) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80143 && (row * 640 + col) <= 80153) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80154 && (row * 640 + col) <= 80181) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80182 && (row * 640 + col) <= 80190) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 80191 && (row * 640 + col) <= 80293) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80294 && (row * 640 + col) <= 80302) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 80303 && (row * 640 + col) <= 80350) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80351 && (row * 640 + col) <= 80357) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80358 && (row * 640 + col) <= 80369) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80370 && (row * 640 + col) <= 80376) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80377 && (row * 640 + col) <= 80486) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80487 && (row * 640 + col) <= 80496) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 80497 && (row * 640 + col) <= 80556) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80557 && (row * 640 + col) <= 80566) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 80567 && (row * 640 + col) <= 80586) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80587 && (row * 640 + col) <= 80595) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80596 && (row * 640 + col) <= 80621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80622 && (row * 640 + col) <= 80629) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80630 && (row * 640 + col) <= 80654) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80655 && (row * 640 + col) <= 80664) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80665 && (row * 640 + col) <= 80782) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80783 && (row * 640 + col) <= 80793) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80794 && (row * 640 + col) <= 80821) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80822 && (row * 640 + col) <= 80830) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 80831 && (row * 640 + col) <= 80933) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80934 && (row * 640 + col) <= 80942) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 80943 && (row * 640 + col) <= 80990) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80991 && (row * 640 + col) <= 80998) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80999 && (row * 640 + col) <= 81008) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81009 && (row * 640 + col) <= 81015) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81016 && (row * 640 + col) <= 81126) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81127 && (row * 640 + col) <= 81136) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 81137 && (row * 640 + col) <= 81196) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81197 && (row * 640 + col) <= 81206) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 81207 && (row * 640 + col) <= 81226) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81227 && (row * 640 + col) <= 81235) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81236 && (row * 640 + col) <= 81261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81262 && (row * 640 + col) <= 81269) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81270 && (row * 640 + col) <= 81294) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81295 && (row * 640 + col) <= 81304) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81305 && (row * 640 + col) <= 81422) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81423 && (row * 640 + col) <= 81433) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81434 && (row * 640 + col) <= 81461) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81462 && (row * 640 + col) <= 81469) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 81470 && (row * 640 + col) <= 81573) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81574 && (row * 640 + col) <= 81582) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 81583 && (row * 640 + col) <= 81631) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81632 && (row * 640 + col) <= 81639) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81640 && (row * 640 + col) <= 81647) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81648 && (row * 640 + col) <= 81654) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81655 && (row * 640 + col) <= 81765) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81766 && (row * 640 + col) <= 81775) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 81776 && (row * 640 + col) <= 81837) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81838 && (row * 640 + col) <= 81846) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 81847 && (row * 640 + col) <= 81866) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81867 && (row * 640 + col) <= 81875) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81876 && (row * 640 + col) <= 81901) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81902 && (row * 640 + col) <= 81910) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81911 && (row * 640 + col) <= 81934) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81935 && (row * 640 + col) <= 81944) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81945 && (row * 640 + col) <= 82062) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82063 && (row * 640 + col) <= 82073) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82074 && (row * 640 + col) <= 82101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82102 && (row * 640 + col) <= 82109) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 82110 && (row * 640 + col) <= 82213) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82214 && (row * 640 + col) <= 82222) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 82223 && (row * 640 + col) <= 82272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82273 && (row * 640 + col) <= 82280) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82281 && (row * 640 + col) <= 82286) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82287 && (row * 640 + col) <= 82293) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82294 && (row * 640 + col) <= 82405) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82406 && (row * 640 + col) <= 82415) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 82416 && (row * 640 + col) <= 82477) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82478 && (row * 640 + col) <= 82487) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 82488 && (row * 640 + col) <= 82507) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82508 && (row * 640 + col) <= 82515) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82516 && (row * 640 + col) <= 82541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82542 && (row * 640 + col) <= 82550) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82551 && (row * 640 + col) <= 82574) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82575 && (row * 640 + col) <= 82584) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82585 && (row * 640 + col) <= 82702) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82703 && (row * 640 + col) <= 82713) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82714 && (row * 640 + col) <= 82741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82742 && (row * 640 + col) <= 82750) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 82751 && (row * 640 + col) <= 82853) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82854 && (row * 640 + col) <= 82862) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 82863 && (row * 640 + col) <= 82885) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82886 && (row * 640 + col) <= 82904) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82905 && (row * 640 + col) <= 82913) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82914 && (row * 640 + col) <= 82921) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82922 && (row * 640 + col) <= 82925) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82926 && (row * 640 + col) <= 82932) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82933 && (row * 640 + col) <= 82941) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82942 && (row * 640 + col) <= 82960) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82961 && (row * 640 + col) <= 83045) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83046 && (row * 640 + col) <= 83055) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 83056 && (row * 640 + col) <= 83117) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83118 && (row * 640 + col) <= 83127) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 83128 && (row * 640 + col) <= 83147) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83148 && (row * 640 + col) <= 83156) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83157 && (row * 640 + col) <= 83181) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83182 && (row * 640 + col) <= 83190) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83191 && (row * 640 + col) <= 83214) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83215 && (row * 640 + col) <= 83224) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83225 && (row * 640 + col) <= 83342) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83343 && (row * 640 + col) <= 83352) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83353 && (row * 640 + col) <= 83381) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83382 && (row * 640 + col) <= 83390) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 83391 && (row * 640 + col) <= 83493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83494 && (row * 640 + col) <= 83502) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 83503 && (row * 640 + col) <= 83523) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83524 && (row * 640 + col) <= 83546) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83547 && (row * 640 + col) <= 83554) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83555 && (row * 640 + col) <= 83571) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83572 && (row * 640 + col) <= 83579) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83580 && (row * 640 + col) <= 83602) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83603 && (row * 640 + col) <= 83685) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83686 && (row * 640 + col) <= 83695) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 83696 && (row * 640 + col) <= 83758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83759 && (row * 640 + col) <= 83767) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 83768 && (row * 640 + col) <= 83787) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83788 && (row * 640 + col) <= 83796) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83797 && (row * 640 + col) <= 83821) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83822 && (row * 640 + col) <= 83830) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83831 && (row * 640 + col) <= 83854) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83855 && (row * 640 + col) <= 83865) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83866 && (row * 640 + col) <= 83982) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83983 && (row * 640 + col) <= 83992) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83993 && (row * 640 + col) <= 84021) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84022 && (row * 640 + col) <= 84030) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 84031 && (row * 640 + col) <= 84132) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84133 && (row * 640 + col) <= 84141) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 84142 && (row * 640 + col) <= 84162) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84163 && (row * 640 + col) <= 84188) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84189 && (row * 640 + col) <= 84195) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84196 && (row * 640 + col) <= 84210) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84211 && (row * 640 + col) <= 84218) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84219 && (row * 640 + col) <= 84244) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84245 && (row * 640 + col) <= 84325) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84326 && (row * 640 + col) <= 84334) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 84335 && (row * 640 + col) <= 84398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84399 && (row * 640 + col) <= 84407) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 84408 && (row * 640 + col) <= 84427) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84428 && (row * 640 + col) <= 84436) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84437 && (row * 640 + col) <= 84461) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84462 && (row * 640 + col) <= 84470) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84471 && (row * 640 + col) <= 84494) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84495 && (row * 640 + col) <= 84505) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84506 && (row * 640 + col) <= 84621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84622 && (row * 640 + col) <= 84632) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84633 && (row * 640 + col) <= 84662) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84663 && (row * 640 + col) <= 84671) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 84672 && (row * 640 + col) <= 84772) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84773 && (row * 640 + col) <= 84781) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 84782 && (row * 640 + col) <= 84801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84802 && (row * 640 + col) <= 84829) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84830 && (row * 640 + col) <= 84836) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84837 && (row * 640 + col) <= 84849) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84850 && (row * 640 + col) <= 84857) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84858 && (row * 640 + col) <= 84885) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84886 && (row * 640 + col) <= 84964) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84965 && (row * 640 + col) <= 84974) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 84975 && (row * 640 + col) <= 85038) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85039 && (row * 640 + col) <= 85047) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 85048 && (row * 640 + col) <= 85067) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85068 && (row * 640 + col) <= 85076) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85077 && (row * 640 + col) <= 85101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85102 && (row * 640 + col) <= 85110) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85111 && (row * 640 + col) <= 85135) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85136 && (row * 640 + col) <= 85146) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85147 && (row * 640 + col) <= 85261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85262 && (row * 640 + col) <= 85272) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85273 && (row * 640 + col) <= 85302) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85303 && (row * 640 + col) <= 85311) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 85312 && (row * 640 + col) <= 85412) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85413 && (row * 640 + col) <= 85421) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 85422 && (row * 640 + col) <= 85440) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85441 && (row * 640 + col) <= 85470) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85471 && (row * 640 + col) <= 85477) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85478 && (row * 640 + col) <= 85488) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85489 && (row * 640 + col) <= 85496) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85497 && (row * 640 + col) <= 85525) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85526 && (row * 640 + col) <= 85604) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85605 && (row * 640 + col) <= 85614) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 85615 && (row * 640 + col) <= 85678) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85679 && (row * 640 + col) <= 85688) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 85689 && (row * 640 + col) <= 85707) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85708 && (row * 640 + col) <= 85716) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85717 && (row * 640 + col) <= 85741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85742 && (row * 640 + col) <= 85750) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85751 && (row * 640 + col) <= 85775) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85776 && (row * 640 + col) <= 85786) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85787 && (row * 640 + col) <= 85900) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85901 && (row * 640 + col) <= 85911) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85912 && (row * 640 + col) <= 85942) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85943 && (row * 640 + col) <= 85952) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 85953 && (row * 640 + col) <= 86051) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86052 && (row * 640 + col) <= 86060) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 86061 && (row * 640 + col) <= 86079) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86080 && (row * 640 + col) <= 86111) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86112 && (row * 640 + col) <= 86118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86119 && (row * 640 + col) <= 86127) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86128 && (row * 640 + col) <= 86135) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86136 && (row * 640 + col) <= 86166) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86167 && (row * 640 + col) <= 86244) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86245 && (row * 640 + col) <= 86254) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 86255 && (row * 640 + col) <= 86318) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86319 && (row * 640 + col) <= 86328) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 86329 && (row * 640 + col) <= 86348) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86349 && (row * 640 + col) <= 86357) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86358 && (row * 640 + col) <= 86381) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86382 && (row * 640 + col) <= 86390) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86391 && (row * 640 + col) <= 86416) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86417 && (row * 640 + col) <= 86426) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86427 && (row * 640 + col) <= 86540) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86541 && (row * 640 + col) <= 86551) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86552 && (row * 640 + col) <= 86583) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86584 && (row * 640 + col) <= 86592) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 86593 && (row * 640 + col) <= 86691) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86692 && (row * 640 + col) <= 86700) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 86701 && (row * 640 + col) <= 86719) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86720 && (row * 640 + col) <= 86726) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86727 && (row * 640 + col) <= 86744) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86745 && (row * 640 + col) <= 86752) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86753 && (row * 640 + col) <= 86760) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86761 && (row * 640 + col) <= 86766) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86767 && (row * 640 + col) <= 86774) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86775 && (row * 640 + col) <= 86782) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86783 && (row * 640 + col) <= 86800) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86801 && (row * 640 + col) <= 86806) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86807 && (row * 640 + col) <= 86884) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86885 && (row * 640 + col) <= 86894) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 86895 && (row * 640 + col) <= 86959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86960 && (row * 640 + col) <= 86968) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 86969 && (row * 640 + col) <= 86988) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86989 && (row * 640 + col) <= 86997) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86998 && (row * 640 + col) <= 87021) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87022 && (row * 640 + col) <= 87030) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87031 && (row * 640 + col) <= 87056) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87057 && (row * 640 + col) <= 87067) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87068 && (row * 640 + col) <= 87180) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87181 && (row * 640 + col) <= 87190) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87191 && (row * 640 + col) <= 87223) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87224 && (row * 640 + col) <= 87232) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 87233 && (row * 640 + col) <= 87330) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87331 && (row * 640 + col) <= 87340) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 87341 && (row * 640 + col) <= 87359) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87360 && (row * 640 + col) <= 87365) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87366 && (row * 640 + col) <= 87385) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87386 && (row * 640 + col) <= 87393) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87394 && (row * 640 + col) <= 87413) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87414 && (row * 640 + col) <= 87420) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87421 && (row * 640 + col) <= 87441) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87442 && (row * 640 + col) <= 87447) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87448 && (row * 640 + col) <= 87524) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87525 && (row * 640 + col) <= 87533) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 87534 && (row * 640 + col) <= 87599) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87600 && (row * 640 + col) <= 87608) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 87609 && (row * 640 + col) <= 87628) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87629 && (row * 640 + col) <= 87637) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87638 && (row * 640 + col) <= 87661) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87662 && (row * 640 + col) <= 87670) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87671 && (row * 640 + col) <= 87696) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87697 && (row * 640 + col) <= 87707) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87708 && (row * 640 + col) <= 87819) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87820 && (row * 640 + col) <= 87830) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87831 && (row * 640 + col) <= 87864) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87865 && (row * 640 + col) <= 87873) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 87874 && (row * 640 + col) <= 87970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87971 && (row * 640 + col) <= 87979) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 87980 && (row * 640 + col) <= 87999) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88000 && (row * 640 + col) <= 88004) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88005 && (row * 640 + col) <= 88026) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88027 && (row * 640 + col) <= 88034) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88035 && (row * 640 + col) <= 88052) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88053 && (row * 640 + col) <= 88059) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88060 && (row * 640 + col) <= 88081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88082 && (row * 640 + col) <= 88087) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88088 && (row * 640 + col) <= 88164) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88165 && (row * 640 + col) <= 88173) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 88174 && (row * 640 + col) <= 88239) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88240 && (row * 640 + col) <= 88248) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 88249 && (row * 640 + col) <= 88268) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88269 && (row * 640 + col) <= 88277) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88278 && (row * 640 + col) <= 88301) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88302 && (row * 640 + col) <= 88310) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88311 && (row * 640 + col) <= 88337) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88338 && (row * 640 + col) <= 88348) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88349 && (row * 640 + col) <= 88459) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88460 && (row * 640 + col) <= 88470) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88471 && (row * 640 + col) <= 88504) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88505 && (row * 640 + col) <= 88513) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 88514 && (row * 640 + col) <= 88610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88611 && (row * 640 + col) <= 88619) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 88620 && (row * 640 + col) <= 88638) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88639 && (row * 640 + col) <= 88644) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88645 && (row * 640 + col) <= 88667) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88668 && (row * 640 + col) <= 88674) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88675 && (row * 640 + col) <= 88691) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88692 && (row * 640 + col) <= 88699) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88700 && (row * 640 + col) <= 88722) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88723 && (row * 640 + col) <= 88727) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88728 && (row * 640 + col) <= 88804) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88805 && (row * 640 + col) <= 88813) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 88814 && (row * 640 + col) <= 88879) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88880 && (row * 640 + col) <= 88888) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 88889 && (row * 640 + col) <= 88908) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88909 && (row * 640 + col) <= 88917) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88918 && (row * 640 + col) <= 88941) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88942 && (row * 640 + col) <= 88950) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88951 && (row * 640 + col) <= 88977) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88978 && (row * 640 + col) <= 88988) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88989 && (row * 640 + col) <= 89098) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89099 && (row * 640 + col) <= 89109) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89110 && (row * 640 + col) <= 89144) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89145 && (row * 640 + col) <= 89154) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 89155 && (row * 640 + col) <= 89249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89250 && (row * 640 + col) <= 89258) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 89259 && (row * 640 + col) <= 89278) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89279 && (row * 640 + col) <= 89284) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89285 && (row * 640 + col) <= 89308) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89309 && (row * 640 + col) <= 89315) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89316 && (row * 640 + col) <= 89331) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89332 && (row * 640 + col) <= 89338) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89339 && (row * 640 + col) <= 89362) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89363 && (row * 640 + col) <= 89367) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89368 && (row * 640 + col) <= 89403) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89404 && (row * 640 + col) <= 89411) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 89412 && (row * 640 + col) <= 89444) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89445 && (row * 640 + col) <= 89453) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 89454 && (row * 640 + col) <= 89519) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89520 && (row * 640 + col) <= 89528) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 89529 && (row * 640 + col) <= 89548) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89549 && (row * 640 + col) <= 89557) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89558 && (row * 640 + col) <= 89581) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89582 && (row * 640 + col) <= 89590) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89591 && (row * 640 + col) <= 89618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89619 && (row * 640 + col) <= 89629) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89630 && (row * 640 + col) <= 89738) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89739 && (row * 640 + col) <= 89749) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89750 && (row * 640 + col) <= 89785) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89786 && (row * 640 + col) <= 89794) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 89795 && (row * 640 + col) <= 89889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89890 && (row * 640 + col) <= 89898) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 89899 && (row * 640 + col) <= 89918) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89919 && (row * 640 + col) <= 89924) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89925 && (row * 640 + col) <= 89949) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89950 && (row * 640 + col) <= 89955) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89956 && (row * 640 + col) <= 89970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89971 && (row * 640 + col) <= 89977) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 89978 && (row * 640 + col) <= 90002) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90003 && (row * 640 + col) <= 90007) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90008 && (row * 640 + col) <= 90039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90040 && (row * 640 + col) <= 90055) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 90056 && (row * 640 + col) <= 90084) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90085 && (row * 640 + col) <= 90093) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 90094 && (row * 640 + col) <= 90159) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90160 && (row * 640 + col) <= 90168) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 90169 && (row * 640 + col) <= 90188) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90189 && (row * 640 + col) <= 90197) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90198 && (row * 640 + col) <= 90221) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90222 && (row * 640 + col) <= 90230) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90231 && (row * 640 + col) <= 90258) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90259 && (row * 640 + col) <= 90269) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90270 && (row * 640 + col) <= 90377) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90378 && (row * 640 + col) <= 90388) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90389 && (row * 640 + col) <= 90425) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90426 && (row * 640 + col) <= 90434) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 90435 && (row * 640 + col) <= 90528) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90529 && (row * 640 + col) <= 90537) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 90538 && (row * 640 + col) <= 90558) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90559 && (row * 640 + col) <= 90564) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90565 && (row * 640 + col) <= 90590) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90591 && (row * 640 + col) <= 90596) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90597 && (row * 640 + col) <= 90610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90611 && (row * 640 + col) <= 90616) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90617 && (row * 640 + col) <= 90642) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90643 && (row * 640 + col) <= 90647) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90648 && (row * 640 + col) <= 90677) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90678 && (row * 640 + col) <= 90698) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 90699 && (row * 640 + col) <= 90724) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90725 && (row * 640 + col) <= 90733) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 90734 && (row * 640 + col) <= 90799) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90800 && (row * 640 + col) <= 90808) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 90809 && (row * 640 + col) <= 90828) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90829 && (row * 640 + col) <= 90837) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90838 && (row * 640 + col) <= 90861) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90862 && (row * 640 + col) <= 90870) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90871 && (row * 640 + col) <= 90898) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90899 && (row * 640 + col) <= 90909) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 90910 && (row * 640 + col) <= 91017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91018 && (row * 640 + col) <= 91028) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91029 && (row * 640 + col) <= 91065) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91066 && (row * 640 + col) <= 91075) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 91076 && (row * 640 + col) <= 91168) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91169 && (row * 640 + col) <= 91177) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 91178 && (row * 640 + col) <= 91198) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91199 && (row * 640 + col) <= 91204) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91205 && (row * 640 + col) <= 91230) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91231 && (row * 640 + col) <= 91236) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91237 && (row * 640 + col) <= 91250) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91251 && (row * 640 + col) <= 91256) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91257 && (row * 640 + col) <= 91282) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91283 && (row * 640 + col) <= 91287) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91288 && (row * 640 + col) <= 91315) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91316 && (row * 640 + col) <= 91340) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 91341 && (row * 640 + col) <= 91364) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91365 && (row * 640 + col) <= 91374) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 91375 && (row * 640 + col) <= 91438) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91439 && (row * 640 + col) <= 91448) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 91449 && (row * 640 + col) <= 91468) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91469 && (row * 640 + col) <= 91477) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91478 && (row * 640 + col) <= 91501) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91502 && (row * 640 + col) <= 91510) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91511 && (row * 640 + col) <= 91539) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91540 && (row * 640 + col) <= 91550) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91551 && (row * 640 + col) <= 91657) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91658 && (row * 640 + col) <= 91667) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91668 && (row * 640 + col) <= 91706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91707 && (row * 640 + col) <= 91715) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 91716 && (row * 640 + col) <= 91807) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91808 && (row * 640 + col) <= 91817) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 91818 && (row * 640 + col) <= 91838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91839 && (row * 640 + col) <= 91844) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91845 && (row * 640 + col) <= 91870) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91871 && (row * 640 + col) <= 91876) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91877 && (row * 640 + col) <= 91890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91891 && (row * 640 + col) <= 91896) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91897 && (row * 640 + col) <= 91922) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91923 && (row * 640 + col) <= 91927) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 91928 && (row * 640 + col) <= 91953) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91954 && (row * 640 + col) <= 91982) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 91983 && (row * 640 + col) <= 92004) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92005 && (row * 640 + col) <= 92014) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 92015 && (row * 640 + col) <= 92078) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92079 && (row * 640 + col) <= 92088) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 92089 && (row * 640 + col) <= 92108) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92109 && (row * 640 + col) <= 92117) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92118 && (row * 640 + col) <= 92141) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92142 && (row * 640 + col) <= 92150) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92151 && (row * 640 + col) <= 92179) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92180 && (row * 640 + col) <= 92190) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92191 && (row * 640 + col) <= 92296) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92297 && (row * 640 + col) <= 92307) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92308 && (row * 640 + col) <= 92346) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92347 && (row * 640 + col) <= 92356) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 92357 && (row * 640 + col) <= 92447) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92448 && (row * 640 + col) <= 92456) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 92457 && (row * 640 + col) <= 92478) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92479 && (row * 640 + col) <= 92484) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92485 && (row * 640 + col) <= 92510) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92511 && (row * 640 + col) <= 92516) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92517 && (row * 640 + col) <= 92530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92531 && (row * 640 + col) <= 92536) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92537 && (row * 640 + col) <= 92562) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92563 && (row * 640 + col) <= 92567) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92568 && (row * 640 + col) <= 92592) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92593 && (row * 640 + col) <= 92623) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 92624 && (row * 640 + col) <= 92644) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92645 && (row * 640 + col) <= 92654) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 92655 && (row * 640 + col) <= 92718) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92719 && (row * 640 + col) <= 92728) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 92729 && (row * 640 + col) <= 92748) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92749 && (row * 640 + col) <= 92756) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92757 && (row * 640 + col) <= 92781) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92782 && (row * 640 + col) <= 92790) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92791 && (row * 640 + col) <= 92820) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92821 && (row * 640 + col) <= 92831) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92832 && (row * 640 + col) <= 92936) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92937 && (row * 640 + col) <= 92947) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 92948 && (row * 640 + col) <= 92987) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92988 && (row * 640 + col) <= 92996) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 92997 && (row * 640 + col) <= 93087) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93088 && (row * 640 + col) <= 93096) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 93097 && (row * 640 + col) <= 93118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93119 && (row * 640 + col) <= 93124) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93125 && (row * 640 + col) <= 93149) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93150 && (row * 640 + col) <= 93155) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93156 && (row * 640 + col) <= 93170) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93171 && (row * 640 + col) <= 93177) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93178 && (row * 640 + col) <= 93202) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93203 && (row * 640 + col) <= 93207) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93208 && (row * 640 + col) <= 93230) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93231 && (row * 640 + col) <= 93265) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 93266 && (row * 640 + col) <= 93285) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93286 && (row * 640 + col) <= 93294) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 93295 && (row * 640 + col) <= 93358) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93359 && (row * 640 + col) <= 93367) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 93368 && (row * 640 + col) <= 93388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93389 && (row * 640 + col) <= 93396) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93397 && (row * 640 + col) <= 93421) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93422 && (row * 640 + col) <= 93430) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93431 && (row * 640 + col) <= 93460) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93461 && (row * 640 + col) <= 93471) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93472 && (row * 640 + col) <= 93576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93577 && (row * 640 + col) <= 93586) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93587 && (row * 640 + col) <= 93627) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93628 && (row * 640 + col) <= 93637) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 93638 && (row * 640 + col) <= 93726) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93727 && (row * 640 + col) <= 93735) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 93736 && (row * 640 + col) <= 93758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93759 && (row * 640 + col) <= 93764) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93765 && (row * 640 + col) <= 93788) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93789 && (row * 640 + col) <= 93795) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93796 && (row * 640 + col) <= 93811) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93812 && (row * 640 + col) <= 93818) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93819 && (row * 640 + col) <= 93842) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93843 && (row * 640 + col) <= 93847) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93848 && (row * 640 + col) <= 93869) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93870 && (row * 640 + col) <= 93906) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 93907 && (row * 640 + col) <= 93925) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93926 && (row * 640 + col) <= 93934) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 93935 && (row * 640 + col) <= 93998) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 93999 && (row * 640 + col) <= 94007) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 94008 && (row * 640 + col) <= 94027) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94028 && (row * 640 + col) <= 94036) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94037 && (row * 640 + col) <= 94061) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94062 && (row * 640 + col) <= 94070) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94071 && (row * 640 + col) <= 94101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94102 && (row * 640 + col) <= 94112) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94113 && (row * 640 + col) <= 94215) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94216 && (row * 640 + col) <= 94226) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94227 && (row * 640 + col) <= 94267) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94268 && (row * 640 + col) <= 94277) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 94278 && (row * 640 + col) <= 94366) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94367 && (row * 640 + col) <= 94375) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 94376 && (row * 640 + col) <= 94398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94399 && (row * 640 + col) <= 94404) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94405 && (row * 640 + col) <= 94427) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94428 && (row * 640 + col) <= 94434) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94435 && (row * 640 + col) <= 94451) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94452 && (row * 640 + col) <= 94459) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94460 && (row * 640 + col) <= 94482) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94483 && (row * 640 + col) <= 94487) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94488 && (row * 640 + col) <= 94508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94509 && (row * 640 + col) <= 94547) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 94548 && (row * 640 + col) <= 94565) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94566 && (row * 640 + col) <= 94575) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 94576 && (row * 640 + col) <= 94638) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94639 && (row * 640 + col) <= 94647) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 94648 && (row * 640 + col) <= 94667) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94668 && (row * 640 + col) <= 94676) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94677 && (row * 640 + col) <= 94701) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94702 && (row * 640 + col) <= 94709) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94710 && (row * 640 + col) <= 94741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94742 && (row * 640 + col) <= 94752) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94753 && (row * 640 + col) <= 94855) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94856 && (row * 640 + col) <= 94865) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94866 && (row * 640 + col) <= 94908) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 94909 && (row * 640 + col) <= 94917) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 94918 && (row * 640 + col) <= 95005) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95006 && (row * 640 + col) <= 95015) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 95016 && (row * 640 + col) <= 95039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95040 && (row * 640 + col) <= 95044) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95045 && (row * 640 + col) <= 95066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95067 && (row * 640 + col) <= 95073) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95074 && (row * 640 + col) <= 95092) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95093 && (row * 640 + col) <= 95100) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95101 && (row * 640 + col) <= 95121) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95122 && (row * 640 + col) <= 95127) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95128 && (row * 640 + col) <= 95147) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95148 && (row * 640 + col) <= 95162) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 95163 && (row * 640 + col) <= 95173) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95174 && (row * 640 + col) <= 95188) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 95189 && (row * 640 + col) <= 95205) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95206 && (row * 640 + col) <= 95215) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 95216 && (row * 640 + col) <= 95277) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95278 && (row * 640 + col) <= 95287) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 95288 && (row * 640 + col) <= 95307) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95308 && (row * 640 + col) <= 95316) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95317 && (row * 640 + col) <= 95341) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95342 && (row * 640 + col) <= 95349) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95350 && (row * 640 + col) <= 95381) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95382 && (row * 640 + col) <= 95392) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95393 && (row * 640 + col) <= 95494) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95495 && (row * 640 + col) <= 95505) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95506 && (row * 640 + col) <= 95548) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95549 && (row * 640 + col) <= 95558) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 95559 && (row * 640 + col) <= 95645) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95646 && (row * 640 + col) <= 95654) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 95655 && (row * 640 + col) <= 95679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95680 && (row * 640 + col) <= 95685) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95686 && (row * 640 + col) <= 95705) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95706 && (row * 640 + col) <= 95713) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95714 && (row * 640 + col) <= 95733) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95734 && (row * 640 + col) <= 95741) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95742 && (row * 640 + col) <= 95761) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95762 && (row * 640 + col) <= 95767) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95768 && (row * 640 + col) <= 95786) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95787 && (row * 640 + col) <= 95799) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 95800 && (row * 640 + col) <= 95816) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95817 && (row * 640 + col) <= 95828) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 95829 && (row * 640 + col) <= 95845) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95846 && (row * 640 + col) <= 95855) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 95856 && (row * 640 + col) <= 95917) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95918 && (row * 640 + col) <= 95926) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 95927 && (row * 640 + col) <= 95947) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95948 && (row * 640 + col) <= 95956) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95957 && (row * 640 + col) <= 95981) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 95982 && (row * 640 + col) <= 95989) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95990 && (row * 640 + col) <= 96022) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96023 && (row * 640 + col) <= 96033) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96034 && (row * 640 + col) <= 96134) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96135 && (row * 640 + col) <= 96145) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96146 && (row * 640 + col) <= 96189) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96190 && (row * 640 + col) <= 96198) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 96199 && (row * 640 + col) <= 96285) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96286 && (row * 640 + col) <= 96294) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 96295 && (row * 640 + col) <= 96319) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96320 && (row * 640 + col) <= 96326) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96327 && (row * 640 + col) <= 96344) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96345 && (row * 640 + col) <= 96352) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96353 && (row * 640 + col) <= 96360) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96361 && (row * 640 + col) <= 96366) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96367 && (row * 640 + col) <= 96374) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96375 && (row * 640 + col) <= 96382) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96383 && (row * 640 + col) <= 96400) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96401 && (row * 640 + col) <= 96406) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96407 && (row * 640 + col) <= 96425) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96426 && (row * 640 + col) <= 96437) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 96438 && (row * 640 + col) <= 96457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96458 && (row * 640 + col) <= 96469) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 96470 && (row * 640 + col) <= 96486) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96487 && (row * 640 + col) <= 96495) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 96496 && (row * 640 + col) <= 96556) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96557 && (row * 640 + col) <= 96566) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 96567 && (row * 640 + col) <= 96587) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96588 && (row * 640 + col) <= 96596) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96597 && (row * 640 + col) <= 96620) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96621 && (row * 640 + col) <= 96629) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96630 && (row * 640 + col) <= 96662) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96663 && (row * 640 + col) <= 96673) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96674 && (row * 640 + col) <= 96774) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96775 && (row * 640 + col) <= 96784) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96785 && (row * 640 + col) <= 96829) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96830 && (row * 640 + col) <= 96839) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 96840 && (row * 640 + col) <= 96924) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96925 && (row * 640 + col) <= 96933) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 96934 && (row * 640 + col) <= 96959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96960 && (row * 640 + col) <= 96991) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96992 && (row * 640 + col) <= 96998) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 96999 && (row * 640 + col) <= 97007) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97008 && (row * 640 + col) <= 97015) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97016 && (row * 640 + col) <= 97046) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97047 && (row * 640 + col) <= 97065) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97066 && (row * 640 + col) <= 97076) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 97077 && (row * 640 + col) <= 97099) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97100 && (row * 640 + col) <= 97110) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 97111 && (row * 640 + col) <= 97126) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97127 && (row * 640 + col) <= 97136) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 97137 && (row * 640 + col) <= 97196) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97197 && (row * 640 + col) <= 97206) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 97207 && (row * 640 + col) <= 97227) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97228 && (row * 640 + col) <= 97236) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97237 && (row * 640 + col) <= 97260) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97261 && (row * 640 + col) <= 97269) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97270 && (row * 640 + col) <= 97303) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97304 && (row * 640 + col) <= 97314) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97315 && (row * 640 + col) <= 97413) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97414 && (row * 640 + col) <= 97424) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97425 && (row * 640 + col) <= 97470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97471 && (row * 640 + col) <= 97479) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 97480 && (row * 640 + col) <= 97564) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97565 && (row * 640 + col) <= 97573) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 97574 && (row * 640 + col) <= 97600) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97601 && (row * 640 + col) <= 97630) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97631 && (row * 640 + col) <= 97637) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97638 && (row * 640 + col) <= 97649) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97650 && (row * 640 + col) <= 97656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97657 && (row * 640 + col) <= 97685) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97686 && (row * 640 + col) <= 97704) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97705 && (row * 640 + col) <= 97715) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 97716 && (row * 640 + col) <= 97740) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97741 && (row * 640 + col) <= 97751) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 97752 && (row * 640 + col) <= 97766) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97767 && (row * 640 + col) <= 97776) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 97777 && (row * 640 + col) <= 97836) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97837 && (row * 640 + col) <= 97846) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 97847 && (row * 640 + col) <= 97867) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97868 && (row * 640 + col) <= 97876) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97877 && (row * 640 + col) <= 97900) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97901 && (row * 640 + col) <= 97909) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97910 && (row * 640 + col) <= 97943) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 97944 && (row * 640 + col) <= 97954) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97955 && (row * 640 + col) <= 98053) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98054 && (row * 640 + col) <= 98063) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98064 && (row * 640 + col) <= 98110) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98111 && (row * 640 + col) <= 98119) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 98120 && (row * 640 + col) <= 98203) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98204 && (row * 640 + col) <= 98212) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 98213 && (row * 640 + col) <= 98241) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98242 && (row * 640 + col) <= 98269) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98270 && (row * 640 + col) <= 98276) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98277 && (row * 640 + col) <= 98290) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98291 && (row * 640 + col) <= 98297) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98298 && (row * 640 + col) <= 98325) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98326 && (row * 640 + col) <= 98344) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98345 && (row * 640 + col) <= 98354) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 98355 && (row * 640 + col) <= 98381) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98382 && (row * 640 + col) <= 98391) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 98392 && (row * 640 + col) <= 98407) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98408 && (row * 640 + col) <= 98417) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 98418 && (row * 640 + col) <= 98475) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98476 && (row * 640 + col) <= 98485) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 98486 && (row * 640 + col) <= 98507) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98508 && (row * 640 + col) <= 98516) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98517 && (row * 640 + col) <= 98539) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98540 && (row * 640 + col) <= 98548) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98549 && (row * 640 + col) <= 98584) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98585 && (row * 640 + col) <= 98594) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98595 && (row * 640 + col) <= 98692) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98693 && (row * 640 + col) <= 98703) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98704 && (row * 640 + col) <= 98750) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98751 && (row * 640 + col) <= 98760) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 98761 && (row * 640 + col) <= 98843) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98844 && (row * 640 + col) <= 98852) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 98853 && (row * 640 + col) <= 98882) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98883 && (row * 640 + col) <= 98908) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98909 && (row * 640 + col) <= 98915) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98916 && (row * 640 + col) <= 98931) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98932 && (row * 640 + col) <= 98938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98939 && (row * 640 + col) <= 98964) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98965 && (row * 640 + col) <= 98983) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 98984 && (row * 640 + col) <= 98993) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 98994 && (row * 640 + col) <= 99022) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99023 && (row * 640 + col) <= 99031) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 99032 && (row * 640 + col) <= 99047) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99048 && (row * 640 + col) <= 99057) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 99058 && (row * 640 + col) <= 99115) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99116 && (row * 640 + col) <= 99125) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 99126 && (row * 640 + col) <= 99147) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99148 && (row * 640 + col) <= 99156) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99157 && (row * 640 + col) <= 99179) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99180 && (row * 640 + col) <= 99188) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99189 && (row * 640 + col) <= 99224) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99225 && (row * 640 + col) <= 99235) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99236 && (row * 640 + col) <= 99332) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99333 && (row * 640 + col) <= 99342) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99343 && (row * 640 + col) <= 99391) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99392 && (row * 640 + col) <= 99400) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 99401 && (row * 640 + col) <= 99482) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99483 && (row * 640 + col) <= 99492) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 99493 && (row * 640 + col) <= 99523) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99524 && (row * 640 + col) <= 99546) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99547 && (row * 640 + col) <= 99554) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99555 && (row * 640 + col) <= 99572) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99573 && (row * 640 + col) <= 99579) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99580 && (row * 640 + col) <= 99602) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99603 && (row * 640 + col) <= 99623) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99624 && (row * 640 + col) <= 99632) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 99633 && (row * 640 + col) <= 99663) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99664 && (row * 640 + col) <= 99672) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 99673 && (row * 640 + col) <= 99687) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99688 && (row * 640 + col) <= 99698) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 99699 && (row * 640 + col) <= 99754) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99755 && (row * 640 + col) <= 99764) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 99765 && (row * 640 + col) <= 99787) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99788 && (row * 640 + col) <= 99796) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99797 && (row * 640 + col) <= 99819) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99820 && (row * 640 + col) <= 99828) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99829 && (row * 640 + col) <= 99864) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99865 && (row * 640 + col) <= 99875) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99876 && (row * 640 + col) <= 99971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 99972 && (row * 640 + col) <= 99982) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99983 && (row * 640 + col) <= 100031) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100032 && (row * 640 + col) <= 100041) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 100042 && (row * 640 + col) <= 100122) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100123 && (row * 640 + col) <= 100131) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 100132 && (row * 640 + col) <= 100165) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100166 && (row * 640 + col) <= 100184) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100185 && (row * 640 + col) <= 100193) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100194 && (row * 640 + col) <= 100201) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100202 && (row * 640 + col) <= 100205) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100206 && (row * 640 + col) <= 100213) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100214 && (row * 640 + col) <= 100221) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100222 && (row * 640 + col) <= 100240) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100241 && (row * 640 + col) <= 100262) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100263 && (row * 640 + col) <= 100271) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 100272 && (row * 640 + col) <= 100303) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100304 && (row * 640 + col) <= 100312) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 100313 && (row * 640 + col) <= 100328) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100329 && (row * 640 + col) <= 100339) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 100340 && (row * 640 + col) <= 100393) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100394 && (row * 640 + col) <= 100404) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 100405 && (row * 640 + col) <= 100427) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100428 && (row * 640 + col) <= 100436) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100437 && (row * 640 + col) <= 100459) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100460 && (row * 640 + col) <= 100468) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100469 && (row * 640 + col) <= 100505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100506 && (row * 640 + col) <= 100516) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100517 && (row * 640 + col) <= 100611) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100612 && (row * 640 + col) <= 100622) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100623 && (row * 640 + col) <= 100672) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100673 && (row * 640 + col) <= 100681) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 100682 && (row * 640 + col) <= 100762) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100763 && (row * 640 + col) <= 100771) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 100772 && (row * 640 + col) <= 100832) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100833 && (row * 640 + col) <= 100840) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100841 && (row * 640 + col) <= 100846) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100847 && (row * 640 + col) <= 100854) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100855 && (row * 640 + col) <= 100902) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100903 && (row * 640 + col) <= 100911) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 100912 && (row * 640 + col) <= 100944) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100945 && (row * 640 + col) <= 100953) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 100954 && (row * 640 + col) <= 100968) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 100969 && (row * 640 + col) <= 100979) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 100980 && (row * 640 + col) <= 101033) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101034 && (row * 640 + col) <= 101043) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 101044 && (row * 640 + col) <= 101067) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101068 && (row * 640 + col) <= 101076) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101077 && (row * 640 + col) <= 101098) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101099 && (row * 640 + col) <= 101107) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101108 && (row * 640 + col) <= 101145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101146 && (row * 640 + col) <= 101156) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101157 && (row * 640 + col) <= 101251) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101252 && (row * 640 + col) <= 101261) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101262 && (row * 640 + col) <= 101312) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101313 && (row * 640 + col) <= 101321) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 101322 && (row * 640 + col) <= 101401) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101402 && (row * 640 + col) <= 101410) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 101411 && (row * 640 + col) <= 101471) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101472 && (row * 640 + col) <= 101479) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101480 && (row * 640 + col) <= 101487) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101488 && (row * 640 + col) <= 101495) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101496 && (row * 640 + col) <= 101542) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101543 && (row * 640 + col) <= 101550) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 101551 && (row * 640 + col) <= 101584) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101585 && (row * 640 + col) <= 101593) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 101594 && (row * 640 + col) <= 101609) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101610 && (row * 640 + col) <= 101620) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 101621 && (row * 640 + col) <= 101672) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101673 && (row * 640 + col) <= 101683) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 101684 && (row * 640 + col) <= 101707) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101708 && (row * 640 + col) <= 101716) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101717 && (row * 640 + col) <= 101738) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101739 && (row * 640 + col) <= 101747) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101748 && (row * 640 + col) <= 101786) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101787 && (row * 640 + col) <= 101797) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101798 && (row * 640 + col) <= 101890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101891 && (row * 640 + col) <= 101901) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101902 && (row * 640 + col) <= 101952) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 101953 && (row * 640 + col) <= 101962) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 101963 && (row * 640 + col) <= 102041) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102042 && (row * 640 + col) <= 102050) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 102051 && (row * 640 + col) <= 102110) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102111 && (row * 640 + col) <= 102118) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102119 && (row * 640 + col) <= 102128) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102129 && (row * 640 + col) <= 102135) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102136 && (row * 640 + col) <= 102181) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102182 && (row * 640 + col) <= 102190) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 102191 && (row * 640 + col) <= 102225) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102226 && (row * 640 + col) <= 102233) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 102234 && (row * 640 + col) <= 102249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102250 && (row * 640 + col) <= 102261) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 102262 && (row * 640 + col) <= 102311) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102312 && (row * 640 + col) <= 102323) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 102324 && (row * 640 + col) <= 102347) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102348 && (row * 640 + col) <= 102356) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102357 && (row * 640 + col) <= 102377) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102378 && (row * 640 + col) <= 102387) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102388 && (row * 640 + col) <= 102426) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102427 && (row * 640 + col) <= 102437) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102438 && (row * 640 + col) <= 102530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102531 && (row * 640 + col) <= 102540) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102541 && (row * 640 + col) <= 102593) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102594 && (row * 640 + col) <= 102602) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 102603 && (row * 640 + col) <= 102680) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102681 && (row * 640 + col) <= 102690) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 102691 && (row * 640 + col) <= 102750) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102751 && (row * 640 + col) <= 102757) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102758 && (row * 640 + col) <= 102769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102770 && (row * 640 + col) <= 102776) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102777 && (row * 640 + col) <= 102821) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102822 && (row * 640 + col) <= 102829) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 102830 && (row * 640 + col) <= 102865) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102866 && (row * 640 + col) <= 102873) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 102874 && (row * 640 + col) <= 102890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102891 && (row * 640 + col) <= 102902) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 102903 && (row * 640 + col) <= 102951) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102952 && (row * 640 + col) <= 102962) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 102963 && (row * 640 + col) <= 102987) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 102988 && (row * 640 + col) <= 102996) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102997 && (row * 640 + col) <= 103016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103017 && (row * 640 + col) <= 103026) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103027 && (row * 640 + col) <= 103066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103067 && (row * 640 + col) <= 103077) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103078 && (row * 640 + col) <= 103169) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103170 && (row * 640 + col) <= 103180) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103181 && (row * 640 + col) <= 103233) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103234 && (row * 640 + col) <= 103243) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 103244 && (row * 640 + col) <= 103320) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103321 && (row * 640 + col) <= 103329) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 103330 && (row * 640 + col) <= 103389) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103390 && (row * 640 + col) <= 103396) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103397 && (row * 640 + col) <= 103410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103411 && (row * 640 + col) <= 103416) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103417 && (row * 640 + col) <= 103461) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103462 && (row * 640 + col) <= 103469) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 103470 && (row * 640 + col) <= 103505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103506 && (row * 640 + col) <= 103514) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 103515 && (row * 640 + col) <= 103530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103531 && (row * 640 + col) <= 103543) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 103544 && (row * 640 + col) <= 103590) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103591 && (row * 640 + col) <= 103601) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 103602 && (row * 640 + col) <= 103628) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103629 && (row * 640 + col) <= 103637) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103638 && (row * 640 + col) <= 103656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103657 && (row * 640 + col) <= 103666) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103667 && (row * 640 + col) <= 103707) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103708 && (row * 640 + col) <= 103718) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103719 && (row * 640 + col) <= 103809) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103810 && (row * 640 + col) <= 103820) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103821 && (row * 640 + col) <= 103874) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103875 && (row * 640 + col) <= 103883) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 103884 && (row * 640 + col) <= 103960) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 103961 && (row * 640 + col) <= 103969) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 103970 && (row * 640 + col) <= 104029) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104030 && (row * 640 + col) <= 104035) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104036 && (row * 640 + col) <= 104051) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104052 && (row * 640 + col) <= 104057) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104058 && (row * 640 + col) <= 104101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104102 && (row * 640 + col) <= 104109) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 104110 && (row * 640 + col) <= 104146) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104147 && (row * 640 + col) <= 104154) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 104155 && (row * 640 + col) <= 104171) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104172 && (row * 640 + col) <= 104183) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 104184 && (row * 640 + col) <= 104229) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104230 && (row * 640 + col) <= 104241) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 104242 && (row * 640 + col) <= 104268) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104269 && (row * 640 + col) <= 104277) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104278 && (row * 640 + col) <= 104295) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104296 && (row * 640 + col) <= 104305) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104306 && (row * 640 + col) <= 104347) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104348 && (row * 640 + col) <= 104358) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104359 && (row * 640 + col) <= 104449) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104450 && (row * 640 + col) <= 104459) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104460 && (row * 640 + col) <= 104514) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104515 && (row * 640 + col) <= 104524) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 104525 && (row * 640 + col) <= 104599) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104600 && (row * 640 + col) <= 104608) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 104609 && (row * 640 + col) <= 104669) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104670 && (row * 640 + col) <= 104674) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104675 && (row * 640 + col) <= 104691) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104692 && (row * 640 + col) <= 104697) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104698 && (row * 640 + col) <= 104741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104742 && (row * 640 + col) <= 104749) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 104750 && (row * 640 + col) <= 104786) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104787 && (row * 640 + col) <= 104794) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 104795 && (row * 640 + col) <= 104812) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104813 && (row * 640 + col) <= 104825) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 104826 && (row * 640 + col) <= 104868) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104869 && (row * 640 + col) <= 104880) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 104881 && (row * 640 + col) <= 104908) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104909 && (row * 640 + col) <= 104918) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104919 && (row * 640 + col) <= 104934) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104935 && (row * 640 + col) <= 104945) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104946 && (row * 640 + col) <= 104988) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 104989 && (row * 640 + col) <= 104999) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105000 && (row * 640 + col) <= 105088) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105089 && (row * 640 + col) <= 105099) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105100 && (row * 640 + col) <= 105155) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105156 && (row * 640 + col) <= 105164) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 105165 && (row * 640 + col) <= 105239) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105240 && (row * 640 + col) <= 105248) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 105249 && (row * 640 + col) <= 105309) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105310 && (row * 640 + col) <= 105314) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105315 && (row * 640 + col) <= 105331) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105332 && (row * 640 + col) <= 105337) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105338 && (row * 640 + col) <= 105380) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105381 && (row * 640 + col) <= 105389) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 105390 && (row * 640 + col) <= 105426) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105427 && (row * 640 + col) <= 105434) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 105435 && (row * 640 + col) <= 105453) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105454 && (row * 640 + col) <= 105466) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 105467 && (row * 640 + col) <= 105506) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105507 && (row * 640 + col) <= 105519) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 105520 && (row * 640 + col) <= 105548) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105549 && (row * 640 + col) <= 105558) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105559 && (row * 640 + col) <= 105573) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105574 && (row * 640 + col) <= 105584) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105585 && (row * 640 + col) <= 105628) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105629 && (row * 640 + col) <= 105639) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105640 && (row * 640 + col) <= 105728) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105729 && (row * 640 + col) <= 105739) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105740 && (row * 640 + col) <= 105795) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105796 && (row * 640 + col) <= 105805) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 105806 && (row * 640 + col) <= 105877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105878 && (row * 640 + col) <= 105887) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 105888 && (row * 640 + col) <= 105949) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105950 && (row * 640 + col) <= 105954) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105955 && (row * 640 + col) <= 105971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 105972 && (row * 640 + col) <= 105977) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105978 && (row * 640 + col) <= 106020) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106021 && (row * 640 + col) <= 106029) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 106030 && (row * 640 + col) <= 106066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106067 && (row * 640 + col) <= 106074) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 106075 && (row * 640 + col) <= 106094) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106095 && (row * 640 + col) <= 106107) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 106108 && (row * 640 + col) <= 106145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106146 && (row * 640 + col) <= 106158) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 106159 && (row * 640 + col) <= 106189) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106190 && (row * 640 + col) <= 106200) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106201 && (row * 640 + col) <= 106212) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106213 && (row * 640 + col) <= 106223) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106224 && (row * 640 + col) <= 106269) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106270 && (row * 640 + col) <= 106279) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106280 && (row * 640 + col) <= 106367) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106368 && (row * 640 + col) <= 106378) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106379 && (row * 640 + col) <= 106435) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106436 && (row * 640 + col) <= 106447) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 106448 && (row * 640 + col) <= 106515) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106516 && (row * 640 + col) <= 106527) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 106528 && (row * 640 + col) <= 106589) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106590 && (row * 640 + col) <= 106594) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106595 && (row * 640 + col) <= 106611) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106612 && (row * 640 + col) <= 106617) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106618 && (row * 640 + col) <= 106660) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106661 && (row * 640 + col) <= 106669) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 106670 && (row * 640 + col) <= 106706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106707 && (row * 640 + col) <= 106714) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 106715 && (row * 640 + col) <= 106734) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106735 && (row * 640 + col) <= 106749) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 106750 && (row * 640 + col) <= 106783) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106784 && (row * 640 + col) <= 106798) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 106799 && (row * 640 + col) <= 106829) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106830 && (row * 640 + col) <= 106841) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106842 && (row * 640 + col) <= 106850) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106851 && (row * 640 + col) <= 106863) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106864 && (row * 640 + col) <= 106909) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 106910 && (row * 640 + col) <= 106920) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106921 && (row * 640 + col) <= 107007) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107008 && (row * 640 + col) <= 107018) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107019 && (row * 640 + col) <= 107076) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107077 && (row * 640 + col) <= 107090) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 107091 && (row * 640 + col) <= 107153) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107154 && (row * 640 + col) <= 107167) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 107168 && (row * 640 + col) <= 107229) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107230 && (row * 640 + col) <= 107234) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107235 && (row * 640 + col) <= 107251) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107252 && (row * 640 + col) <= 107257) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107258 && (row * 640 + col) <= 107300) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107301 && (row * 640 + col) <= 107309) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 107310 && (row * 640 + col) <= 107346) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107347 && (row * 640 + col) <= 107354) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 107355 && (row * 640 + col) <= 107375) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107376 && (row * 640 + col) <= 107390) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 107391 && (row * 640 + col) <= 107422) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107423 && (row * 640 + col) <= 107437) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 107438 && (row * 640 + col) <= 107470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107471 && (row * 640 + col) <= 107484) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107485 && (row * 640 + col) <= 107487) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107488 && (row * 640 + col) <= 107502) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107503 && (row * 640 + col) <= 107549) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107550 && (row * 640 + col) <= 107560) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107561 && (row * 640 + col) <= 107646) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107647 && (row * 640 + col) <= 107657) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107658 && (row * 640 + col) <= 107716) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107717 && (row * 640 + col) <= 107732) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 107733 && (row * 640 + col) <= 107790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107791 && (row * 640 + col) <= 107806) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 107807 && (row * 640 + col) <= 107869) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107870 && (row * 640 + col) <= 107874) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107875 && (row * 640 + col) <= 107891) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107892 && (row * 640 + col) <= 107897) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107898 && (row * 640 + col) <= 107940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107941 && (row * 640 + col) <= 107949) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 107950 && (row * 640 + col) <= 107986) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 107987 && (row * 640 + col) <= 107994) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 107995 && (row * 640 + col) <= 108016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108017 && (row * 640 + col) <= 108032) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 108033 && (row * 640 + col) <= 108060) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108061 && (row * 640 + col) <= 108076) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 108077 && (row * 640 + col) <= 108110) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108111 && (row * 640 + col) <= 108141) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108142 && (row * 640 + col) <= 108190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108191 && (row * 640 + col) <= 108201) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108202 && (row * 640 + col) <= 108286) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108287 && (row * 640 + col) <= 108297) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108298 && (row * 640 + col) <= 108357) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108358 && (row * 640 + col) <= 108375) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 108376 && (row * 640 + col) <= 108428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108429 && (row * 640 + col) <= 108445) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 108446 && (row * 640 + col) <= 108509) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108510 && (row * 640 + col) <= 108514) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108515 && (row * 640 + col) <= 108531) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108532 && (row * 640 + col) <= 108537) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108538 && (row * 640 + col) <= 108581) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108582 && (row * 640 + col) <= 108589) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 108590 && (row * 640 + col) <= 108626) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108627 && (row * 640 + col) <= 108634) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 108635 && (row * 640 + col) <= 108657) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108658 && (row * 640 + col) <= 108675) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 108676 && (row * 640 + col) <= 108697) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108698 && (row * 640 + col) <= 108715) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 108716 && (row * 640 + col) <= 108751) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108752 && (row * 640 + col) <= 108780) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108781 && (row * 640 + col) <= 108830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108831 && (row * 640 + col) <= 108842) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108843 && (row * 640 + col) <= 108925) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108926 && (row * 640 + col) <= 108936) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108937 && (row * 640 + col) <= 108998) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 108999 && (row * 640 + col) <= 109017) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 109018 && (row * 640 + col) <= 109066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109067 && (row * 640 + col) <= 109085) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 109086 && (row * 640 + col) <= 109149) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109150 && (row * 640 + col) <= 109154) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109155 && (row * 640 + col) <= 109171) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109172 && (row * 640 + col) <= 109177) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109178 && (row * 640 + col) <= 109221) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109222 && (row * 640 + col) <= 109229) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 109230 && (row * 640 + col) <= 109266) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109267 && (row * 640 + col) <= 109274) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 109275 && (row * 640 + col) <= 109299) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109300 && (row * 640 + col) <= 109317) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 109318 && (row * 640 + col) <= 109335) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109336 && (row * 640 + col) <= 109353) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 109354 && (row * 640 + col) <= 109392) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109393 && (row * 640 + col) <= 109419) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109420 && (row * 640 + col) <= 109471) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109472 && (row * 640 + col) <= 109484) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109485 && (row * 640 + col) <= 109563) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109564 && (row * 640 + col) <= 109576) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109577 && (row * 640 + col) <= 109639) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109640 && (row * 640 + col) <= 109660) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 109661 && (row * 640 + col) <= 109703) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109704 && (row * 640 + col) <= 109724) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 109725 && (row * 640 + col) <= 109789) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109790 && (row * 640 + col) <= 109794) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109795 && (row * 640 + col) <= 109811) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109812 && (row * 640 + col) <= 109817) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109818 && (row * 640 + col) <= 109861) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109862 && (row * 640 + col) <= 109869) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 109870 && (row * 640 + col) <= 109905) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109906 && (row * 640 + col) <= 109914) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 109915 && (row * 640 + col) <= 109940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109941 && (row * 640 + col) <= 109963) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 109964 && (row * 640 + col) <= 109969) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 109970 && (row * 640 + col) <= 109992) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 109993 && (row * 640 + col) <= 110033) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110034 && (row * 640 + col) <= 110058) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110059 && (row * 640 + col) <= 110111) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110112 && (row * 640 + col) <= 110126) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110127 && (row * 640 + col) <= 110201) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110202 && (row * 640 + col) <= 110216) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110217 && (row * 640 + col) <= 110280) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110281 && (row * 640 + col) <= 110302) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 110303 && (row * 640 + col) <= 110341) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110342 && (row * 640 + col) <= 110362) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 110363 && (row * 640 + col) <= 110429) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110430 && (row * 640 + col) <= 110434) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110435 && (row * 640 + col) <= 110451) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110452 && (row * 640 + col) <= 110457) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110458 && (row * 640 + col) <= 110501) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110502 && (row * 640 + col) <= 110510) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 110511 && (row * 640 + col) <= 110545) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110546 && (row * 640 + col) <= 110553) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 110554 && (row * 640 + col) <= 110581) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110582 && (row * 640 + col) <= 110631) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 110632 && (row * 640 + col) <= 110674) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110675 && (row * 640 + col) <= 110697) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110698 && (row * 640 + col) <= 110752) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110753 && (row * 640 + col) <= 110769) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110770 && (row * 640 + col) <= 110838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110839 && (row * 640 + col) <= 110855) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110856 && (row * 640 + col) <= 110922) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110923 && (row * 640 + col) <= 110944) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 110945 && (row * 640 + col) <= 110979) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 110980 && (row * 640 + col) <= 111001) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 111002 && (row * 640 + col) <= 111069) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111070 && (row * 640 + col) <= 111074) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111075 && (row * 640 + col) <= 111091) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111092 && (row * 640 + col) <= 111097) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111098 && (row * 640 + col) <= 111141) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111142 && (row * 640 + col) <= 111150) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 111151 && (row * 640 + col) <= 111185) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111186 && (row * 640 + col) <= 111193) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 111194 && (row * 640 + col) <= 111223) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111224 && (row * 640 + col) <= 111269) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 111270 && (row * 640 + col) <= 111316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111317 && (row * 640 + col) <= 111335) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111336 && (row * 640 + col) <= 111392) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111393 && (row * 640 + col) <= 111411) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111412 && (row * 640 + col) <= 111476) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111477 && (row * 640 + col) <= 111494) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111495 && (row * 640 + col) <= 111564) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111565 && (row * 640 + col) <= 111587) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 111588 && (row * 640 + col) <= 111616) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111617 && (row * 640 + col) <= 111638) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 111639 && (row * 640 + col) <= 111709) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111710 && (row * 640 + col) <= 111714) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111715 && (row * 640 + col) <= 111731) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111732 && (row * 640 + col) <= 111737) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111738 && (row * 640 + col) <= 111782) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111783 && (row * 640 + col) <= 111791) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 111792 && (row * 640 + col) <= 111824) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111825 && (row * 640 + col) <= 111833) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 111834 && (row * 640 + col) <= 111864) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111865 && (row * 640 + col) <= 111908) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 111909 && (row * 640 + col) <= 111958) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 111959 && (row * 640 + col) <= 111973) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111974 && (row * 640 + col) <= 112033) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112034 && (row * 640 + col) <= 112053) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112054 && (row * 640 + col) <= 112113) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112114 && (row * 640 + col) <= 112134) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112135 && (row * 640 + col) <= 112207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112208 && (row * 640 + col) <= 112229) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 112230 && (row * 640 + col) <= 112254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112255 && (row * 640 + col) <= 112276) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 112277 && (row * 640 + col) <= 112349) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112350 && (row * 640 + col) <= 112354) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112355 && (row * 640 + col) <= 112371) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112372 && (row * 640 + col) <= 112377) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112378 && (row * 640 + col) <= 112422) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112423 && (row * 640 + col) <= 112431) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 112432 && (row * 640 + col) <= 112464) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112465 && (row * 640 + col) <= 112473) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 112474 && (row * 640 + col) <= 112506) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112507 && (row * 640 + col) <= 112547) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 112548 && (row * 640 + col) <= 112600) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112601 && (row * 640 + col) <= 112611) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112612 && (row * 640 + col) <= 112674) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112675 && (row * 640 + col) <= 112696) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112697 && (row * 640 + col) <= 112751) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112752 && (row * 640 + col) <= 112773) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112774 && (row * 640 + col) <= 112849) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112850 && (row * 640 + col) <= 112872) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 112873 && (row * 640 + col) <= 112891) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112892 && (row * 640 + col) <= 112913) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 112914 && (row * 640 + col) <= 112989) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 112990 && (row * 640 + col) <= 112994) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112995 && (row * 640 + col) <= 113011) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113012 && (row * 640 + col) <= 113017) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 113018 && (row * 640 + col) <= 113062) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113063 && (row * 640 + col) <= 113072) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 113073 && (row * 640 + col) <= 113103) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113104 && (row * 640 + col) <= 113112) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 113113 && (row * 640 + col) <= 113148) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113149 && (row * 640 + col) <= 113184) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 113185 && (row * 640 + col) <= 113315) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113316 && (row * 640 + col) <= 113338) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 113339 && (row * 640 + col) <= 113388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113389 && (row * 640 + col) <= 113412) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 113413 && (row * 640 + col) <= 113491) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113492 && (row * 640 + col) <= 113514) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 113515 && (row * 640 + col) <= 113529) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113530 && (row * 640 + col) <= 113551) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 113552 && (row * 640 + col) <= 113629) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113630 && (row * 640 + col) <= 113634) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 113635 && (row * 640 + col) <= 113651) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113652 && (row * 640 + col) <= 113657) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 113658 && (row * 640 + col) <= 113703) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113704 && (row * 640 + col) <= 113712) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 113713 && (row * 640 + col) <= 113742) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113743 && (row * 640 + col) <= 113752) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 113753 && (row * 640 + col) <= 113790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113791 && (row * 640 + col) <= 113822) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 113823 && (row * 640 + col) <= 113956) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 113957 && (row * 640 + col) <= 113981) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 113982 && (row * 640 + col) <= 114026) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114027 && (row * 640 + col) <= 114051) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114052 && (row * 640 + col) <= 114134) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114135 && (row * 640 + col) <= 114156) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 114157 && (row * 640 + col) <= 114167) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114168 && (row * 640 + col) <= 114189) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 114190 && (row * 640 + col) <= 114269) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114270 && (row * 640 + col) <= 114275) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114276 && (row * 640 + col) <= 114291) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114292 && (row * 640 + col) <= 114296) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114297 && (row * 640 + col) <= 114343) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114344 && (row * 640 + col) <= 114353) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 114354 && (row * 640 + col) <= 114382) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114383 && (row * 640 + col) <= 114391) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 114392 && (row * 640 + col) <= 114433) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114434 && (row * 640 + col) <= 114459) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 114460 && (row * 640 + col) <= 114598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114599 && (row * 640 + col) <= 114623) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114624 && (row * 640 + col) <= 114663) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114664 && (row * 640 + col) <= 114689) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114690 && (row * 640 + col) <= 114776) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114777 && (row * 640 + col) <= 114799) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 114800 && (row * 640 + col) <= 114804) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114805 && (row * 640 + col) <= 114826) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 114827 && (row * 640 + col) <= 114909) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114910 && (row * 640 + col) <= 114915) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114916 && (row * 640 + col) <= 114931) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114932 && (row * 640 + col) <= 114936) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114937 && (row * 640 + col) <= 114984) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 114985 && (row * 640 + col) <= 114994) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 114995 && (row * 640 + col) <= 115021) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115022 && (row * 640 + col) <= 115031) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 115032 && (row * 640 + col) <= 115076) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115077 && (row * 640 + col) <= 115096) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 115097 && (row * 640 + col) <= 115239) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115240 && (row * 640 + col) <= 115265) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115266 && (row * 640 + col) <= 115301) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115302 && (row * 640 + col) <= 115327) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115328 && (row * 640 + col) <= 115419) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115420 && (row * 640 + col) <= 115464) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 115465 && (row * 640 + col) <= 115549) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115550 && (row * 640 + col) <= 115556) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115557 && (row * 640 + col) <= 115570) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115571 && (row * 640 + col) <= 115576) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115577 && (row * 640 + col) <= 115624) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115625 && (row * 640 + col) <= 115635) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 115636 && (row * 640 + col) <= 115660) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115661 && (row * 640 + col) <= 115670) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 115671 && (row * 640 + col) <= 115720) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115721 && (row * 640 + col) <= 115732) color_data <= 12'b011111110111; else
        if ((row * 640 + col) >= 115733 && (row * 640 + col) <= 115882) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115883 && (row * 640 + col) <= 115908) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115909 && (row * 640 + col) <= 115939) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 115940 && (row * 640 + col) <= 115965) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115966 && (row * 640 + col) <= 116061) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116062 && (row * 640 + col) <= 116101) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 116102 && (row * 640 + col) <= 116190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116191 && (row * 640 + col) <= 116197) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 116198 && (row * 640 + col) <= 116208) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116209 && (row * 640 + col) <= 116216) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 116217 && (row * 640 + col) <= 116265) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116266 && (row * 640 + col) <= 116276) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 116277 && (row * 640 + col) <= 116298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116299 && (row * 640 + col) <= 116309) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 116310 && (row * 640 + col) <= 116524) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116525 && (row * 640 + col) <= 116550) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 116551 && (row * 640 + col) <= 116576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116577 && (row * 640 + col) <= 116602) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 116603 && (row * 640 + col) <= 116704) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116705 && (row * 640 + col) <= 116739) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 116740 && (row * 640 + col) <= 116830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116831 && (row * 640 + col) <= 116855) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 116856 && (row * 640 + col) <= 116906) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116907 && (row * 640 + col) <= 116918) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 116919 && (row * 640 + col) <= 116937) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 116938 && (row * 640 + col) <= 116949) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 116950 && (row * 640 + col) <= 117166) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117167 && (row * 640 + col) <= 117193) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 117194 && (row * 640 + col) <= 117214) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117215 && (row * 640 + col) <= 117240) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 117241 && (row * 640 + col) <= 117346) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117347 && (row * 640 + col) <= 117377) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 117378 && (row * 640 + col) <= 117471) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117472 && (row * 640 + col) <= 117494) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 117495 && (row * 640 + col) <= 117547) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117548 && (row * 640 + col) <= 117560) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 117561 && (row * 640 + col) <= 117575) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117576 && (row * 640 + col) <= 117588) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 117589 && (row * 640 + col) <= 117809) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117810 && (row * 640 + col) <= 117835) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 117836 && (row * 640 + col) <= 117851) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117852 && (row * 640 + col) <= 117877) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 117878 && (row * 640 + col) <= 117989) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 117990 && (row * 640 + col) <= 118014) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 118015 && (row * 640 + col) <= 118112) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118113 && (row * 640 + col) <= 118134) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 118135 && (row * 640 + col) <= 118187) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118188 && (row * 640 + col) <= 118202) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 118203 && (row * 640 + col) <= 118213) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118214 && (row * 640 + col) <= 118227) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 118228 && (row * 640 + col) <= 118451) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118452 && (row * 640 + col) <= 118478) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 118479 && (row * 640 + col) <= 118489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118490 && (row * 640 + col) <= 118515) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 118516 && (row * 640 + col) <= 118631) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118632 && (row * 640 + col) <= 118652) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 118653 && (row * 640 + col) <= 118753) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118754 && (row * 640 + col) <= 118773) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 118774 && (row * 640 + col) <= 118828) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 118829 && (row * 640 + col) <= 118866) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 118867 && (row * 640 + col) <= 119094) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 119095 && (row * 640 + col) <= 119120) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119121 && (row * 640 + col) <= 119127) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 119128 && (row * 640 + col) <= 119153) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119154 && (row * 640 + col) <= 119273) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 119274 && (row * 640 + col) <= 119290) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 119291 && (row * 640 + col) <= 119394) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 119395 && (row * 640 + col) <= 119411) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119412 && (row * 640 + col) <= 119469) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 119470 && (row * 640 + col) <= 119505) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 119506 && (row * 640 + col) <= 119736) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 119737 && (row * 640 + col) <= 119790) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119791 && (row * 640 + col) <= 119916) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 119917 && (row * 640 + col) <= 119927) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 119928 && (row * 640 + col) <= 120111) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 120112 && (row * 640 + col) <= 120144) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 120145 && (row * 640 + col) <= 120379) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 120380 && (row * 640 + col) <= 120428) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 120429 && (row * 640 + col) <= 120559) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 120560 && (row * 640 + col) <= 120564) color_data <= 12'b111111100011; else
        if ((row * 640 + col) >= 120565 && (row * 640 + col) <= 120752) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 120753 && (row * 640 + col) <= 120782) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 120783 && (row * 640 + col) <= 121021) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 121022 && (row * 640 + col) <= 121065) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 121066 && (row * 640 + col) <= 121394) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 121395 && (row * 640 + col) <= 121421) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 121422 && (row * 640 + col) <= 121663) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 121664 && (row * 640 + col) <= 121703) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 121704 && (row * 640 + col) <= 122035) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 122036 && (row * 640 + col) <= 122059) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 122060 && (row * 640 + col) <= 122306) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 122307 && (row * 640 + col) <= 122341) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 122342 && (row * 640 + col) <= 122678) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 122679 && (row * 640 + col) <= 122697) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 122698 && (row * 640 + col) <= 122949) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 122950 && (row * 640 + col) <= 122978) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 122979 && (row * 640 + col) <= 123321) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 123322 && (row * 640 + col) <= 123333) color_data <= 12'b111100100101; else
        if ((row * 640 + col) >= 123334 && (row * 640 + col) <= 123591) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 123592 && (row * 640 + col) <= 123616) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 123617 && (row * 640 + col) <= 124233) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 124234 && (row * 640 + col) <= 124254) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 124255 && (row * 640 + col) <= 124876) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 124877 && (row * 640 + col) <= 124891) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 124892 && (row * 640 + col) <= 125518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 125519 && (row * 640 + col) <= 125529) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 125530 && (row * 640 + col) < 142720) color_data <= 12'b000000000000; else
        color_data <= 12'b000000000000;
    end
endmodule
