`timescale 1ns / 1ps
module test_rom (
    input wire clk,
    input wire [7:0] row,
    input wire [9:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 584 + col) >= 0 && (row * 584 + col) <= 1) color_data <= 12'b100000000001; else
        if ((row * 584 + col) >= 2 && (row * 584 + col) <= 583) color_data <= 12'b110010111110; else
        if ((row * 584 + col) >= 584 && (row * 584 + col) <= 585) color_data <= 12'b100000000001; else
        if ((row * 584 + col) >= 586 && (row * 584 + col) <= 44383) color_data <= 12'b110010111110; else
        if ((row * 584 + col) >= 44384 && (row * 584 + col) <= 44600) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 44601 && (row * 584 + col) <= 44967) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 44968 && (row * 584 + col) <= 45184) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 45185 && (row * 584 + col) <= 45551) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 45552 && (row * 584 + col) <= 45768) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 45769 && (row * 584 + col) <= 46135) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 46136 && (row * 584 + col) <= 46352) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 46353 && (row * 584 + col) <= 46719) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 46720 && (row * 584 + col) <= 46936) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 46937 && (row * 584 + col) <= 47200) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 47201 && (row * 584 + col) <= 47209) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 47210 && (row * 584 + col) <= 47303) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 47304 && (row * 584 + col) <= 47520) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 47521 && (row * 584 + col) <= 47779) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 47780 && (row * 584 + col) <= 47798) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 47799 && (row * 584 + col) <= 47887) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 47888 && (row * 584 + col) <= 48104) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 48105 && (row * 584 + col) <= 48360) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 48361 && (row * 584 + col) <= 48385) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 48386 && (row * 584 + col) <= 48471) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 48472 && (row * 584 + col) <= 48688) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 48689 && (row * 584 + col) <= 48942) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 48943 && (row * 584 + col) <= 48971) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 48972 && (row * 584 + col) <= 49055) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 49056 && (row * 584 + col) <= 49272) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 49273 && (row * 584 + col) <= 49524) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 49525 && (row * 584 + col) <= 49557) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 49558 && (row * 584 + col) <= 49639) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 49640 && (row * 584 + col) <= 49856) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 49857 && (row * 584 + col) <= 50106) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 50107 && (row * 584 + col) <= 50143) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 50144 && (row * 584 + col) <= 50223) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 50224 && (row * 584 + col) <= 50440) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 50441 && (row * 584 + col) <= 50689) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 50690 && (row * 584 + col) <= 50728) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 50729 && (row * 584 + col) <= 50807) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 50808 && (row * 584 + col) <= 51024) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 51025 && (row * 584 + col) <= 51272) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 51273 && (row * 584 + col) <= 51313) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 51314 && (row * 584 + col) <= 51391) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 51392 && (row * 584 + col) <= 51608) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 51609 && (row * 584 + col) <= 51855) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 51856 && (row * 584 + col) <= 51898) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 51899 && (row * 584 + col) <= 51975) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 51976 && (row * 584 + col) <= 52192) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 52193 && (row * 584 + col) <= 52438) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 52439 && (row * 584 + col) <= 52483) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 52484 && (row * 584 + col) <= 52559) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 52560 && (row * 584 + col) <= 52776) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 52777 && (row * 584 + col) <= 53021) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 53022 && (row * 584 + col) <= 53068) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 53069 && (row * 584 + col) <= 53143) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 53144 && (row * 584 + col) <= 53360) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 53361 && (row * 584 + col) <= 53604) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 53605 && (row * 584 + col) <= 53653) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 53654 && (row * 584 + col) <= 53727) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 53728 && (row * 584 + col) <= 53944) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 53945 && (row * 584 + col) <= 54187) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 54188 && (row * 584 + col) <= 54238) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 54239 && (row * 584 + col) <= 54311) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 54312 && (row * 584 + col) <= 54528) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 54529 && (row * 584 + col) <= 54770) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 54771 && (row * 584 + col) <= 54823) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 54824 && (row * 584 + col) <= 54895) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 54896 && (row * 584 + col) <= 55112) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 55113 && (row * 584 + col) <= 55353) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 55354 && (row * 584 + col) <= 55408) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 55409 && (row * 584 + col) <= 55479) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 55480 && (row * 584 + col) <= 55696) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 55697 && (row * 584 + col) <= 55937) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 55938 && (row * 584 + col) <= 55992) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 55993 && (row * 584 + col) <= 56063) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 56064 && (row * 584 + col) <= 56280) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 56281 && (row * 584 + col) <= 56520) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 56521 && (row * 584 + col) <= 56577) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 56578 && (row * 584 + col) <= 56647) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 56648 && (row * 584 + col) <= 56864) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 56865 && (row * 584 + col) <= 57104) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 57105 && (row * 584 + col) <= 57161) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 57162 && (row * 584 + col) <= 57231) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 57232 && (row * 584 + col) <= 57448) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 57449 && (row * 584 + col) <= 57687) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 57688 && (row * 584 + col) <= 57746) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 57747 && (row * 584 + col) <= 57815) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 57816 && (row * 584 + col) <= 58032) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 58033 && (row * 584 + col) <= 58271) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 58272 && (row * 584 + col) <= 58330) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 58331 && (row * 584 + col) <= 58399) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 58400 && (row * 584 + col) <= 58616) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 58617 && (row * 584 + col) <= 58854) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 58855 && (row * 584 + col) <= 58915) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 58916 && (row * 584 + col) <= 58983) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 58984 && (row * 584 + col) <= 59200) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 59201 && (row * 584 + col) <= 59438) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 59439 && (row * 584 + col) <= 59499) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 59500 && (row * 584 + col) <= 59567) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 59568 && (row * 584 + col) <= 59784) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 59785 && (row * 584 + col) <= 60022) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 60023 && (row * 584 + col) <= 60083) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 60084 && (row * 584 + col) <= 60151) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 60152 && (row * 584 + col) <= 60368) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 60369 && (row * 584 + col) <= 60605) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 60606 && (row * 584 + col) <= 60668) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 60669 && (row * 584 + col) <= 60735) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 60736 && (row * 584 + col) <= 60952) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 60953 && (row * 584 + col) <= 61189) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 61190 && (row * 584 + col) <= 61252) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 61253 && (row * 584 + col) <= 61319) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 61320 && (row * 584 + col) <= 61536) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 61537 && (row * 584 + col) <= 61773) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 61774 && (row * 584 + col) <= 61836) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 61837 && (row * 584 + col) <= 61903) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 61904 && (row * 584 + col) <= 62120) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 62121 && (row * 584 + col) <= 62357) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 62358 && (row * 584 + col) <= 62420) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 62421 && (row * 584 + col) <= 62487) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 62488 && (row * 584 + col) <= 62704) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 62705 && (row * 584 + col) <= 62941) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 62942 && (row * 584 + col) <= 63005) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 63006 && (row * 584 + col) <= 63071) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 63072 && (row * 584 + col) <= 63288) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 63289 && (row * 584 + col) <= 63524) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 63525 && (row * 584 + col) <= 63589) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 63590 && (row * 584 + col) <= 63655) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 63656 && (row * 584 + col) <= 63872) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 63873 && (row * 584 + col) <= 64108) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 64109 && (row * 584 + col) <= 64173) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 64174 && (row * 584 + col) <= 64239) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 64240 && (row * 584 + col) <= 64456) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 64457 && (row * 584 + col) <= 64692) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 64693 && (row * 584 + col) <= 64757) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 64758 && (row * 584 + col) <= 64823) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 64824 && (row * 584 + col) <= 65040) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 65041 && (row * 584 + col) <= 65276) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 65277 && (row * 584 + col) <= 65341) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 65342 && (row * 584 + col) <= 65407) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 65408 && (row * 584 + col) <= 65624) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 65625 && (row * 584 + col) <= 65860) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 65861 && (row * 584 + col) <= 65925) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 65926 && (row * 584 + col) <= 65991) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 65992 && (row * 584 + col) <= 66208) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 66209 && (row * 584 + col) <= 66444) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 66445 && (row * 584 + col) <= 66509) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 66510 && (row * 584 + col) <= 66575) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 66576 && (row * 584 + col) <= 66792) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 66793 && (row * 584 + col) <= 67028) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 67029 && (row * 584 + col) <= 67093) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 67094 && (row * 584 + col) <= 67159) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 67160 && (row * 584 + col) <= 67376) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 67377 && (row * 584 + col) <= 67612) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 67613 && (row * 584 + col) <= 67677) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 67678 && (row * 584 + col) <= 67743) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 67744 && (row * 584 + col) <= 67960) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 67961 && (row * 584 + col) <= 68196) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 68197 && (row * 584 + col) <= 68261) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 68262 && (row * 584 + col) <= 68327) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 68328 && (row * 584 + col) <= 68544) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 68545 && (row * 584 + col) <= 68781) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 68782 && (row * 584 + col) <= 68845) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 68846 && (row * 584 + col) <= 68911) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 68912 && (row * 584 + col) <= 69128) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 69129 && (row * 584 + col) <= 69365) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 69366 && (row * 584 + col) <= 69428) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 69429 && (row * 584 + col) <= 69495) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 69496 && (row * 584 + col) <= 69712) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 69713 && (row * 584 + col) <= 69949) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 69950 && (row * 584 + col) <= 70012) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 70013 && (row * 584 + col) <= 70079) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 70080 && (row * 584 + col) <= 70296) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 70297 && (row * 584 + col) <= 70533) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 70534 && (row * 584 + col) <= 70596) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 70597 && (row * 584 + col) <= 70663) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 70664 && (row * 584 + col) <= 70880) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 70881 && (row * 584 + col) <= 71117) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 71118 && (row * 584 + col) <= 71180) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 71181 && (row * 584 + col) <= 71247) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 71248 && (row * 584 + col) <= 71464) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 71465 && (row * 584 + col) <= 71702) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 71703 && (row * 584 + col) <= 71763) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 71764 && (row * 584 + col) <= 71831) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 71832 && (row * 584 + col) <= 72048) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 72049 && (row * 584 + col) <= 72286) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 72287 && (row * 584 + col) <= 72347) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 72348 && (row * 584 + col) <= 72415) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 72416 && (row * 584 + col) <= 72632) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 72633 && (row * 584 + col) <= 72870) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 72871 && (row * 584 + col) <= 72931) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 72932 && (row * 584 + col) <= 72999) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 73000 && (row * 584 + col) <= 73216) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 73217 && (row * 584 + col) <= 73455) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 73456 && (row * 584 + col) <= 73514) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 73515 && (row * 584 + col) <= 73583) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 73584 && (row * 584 + col) <= 73800) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 73801 && (row * 584 + col) <= 74039) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 74040 && (row * 584 + col) <= 74098) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 74099 && (row * 584 + col) <= 74167) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 74168 && (row * 584 + col) <= 74384) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 74385 && (row * 584 + col) <= 74624) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 74625 && (row * 584 + col) <= 74681) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 74682 && (row * 584 + col) <= 74751) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 74752 && (row * 584 + col) <= 74968) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 74969 && (row * 584 + col) <= 75208) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 75209 && (row * 584 + col) <= 75265) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 75266 && (row * 584 + col) <= 75335) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 75336 && (row * 584 + col) <= 75552) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 75553 && (row * 584 + col) <= 75793) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 75794 && (row * 584 + col) <= 75848) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 75849 && (row * 584 + col) <= 75919) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 75920 && (row * 584 + col) <= 76136) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 76137 && (row * 584 + col) <= 76377) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 76378 && (row * 584 + col) <= 76432) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 76433 && (row * 584 + col) <= 76503) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 76504 && (row * 584 + col) <= 76720) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 76721 && (row * 584 + col) <= 76962) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 76963 && (row * 584 + col) <= 77015) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 77016 && (row * 584 + col) <= 77087) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 77088 && (row * 584 + col) <= 77304) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 77305 && (row * 584 + col) <= 77547) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 77548 && (row * 584 + col) <= 77598) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 77599 && (row * 584 + col) <= 77671) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 77672 && (row * 584 + col) <= 77888) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 77889 && (row * 584 + col) <= 78132) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 78133 && (row * 584 + col) <= 78181) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 78182 && (row * 584 + col) <= 78255) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 78256 && (row * 584 + col) <= 78472) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 78473 && (row * 584 + col) <= 78717) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 78718 && (row * 584 + col) <= 78764) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 78765 && (row * 584 + col) <= 78839) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 78840 && (row * 584 + col) <= 79056) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 79057 && (row * 584 + col) <= 79302) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 79303 && (row * 584 + col) <= 79348) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 79349 && (row * 584 + col) <= 79423) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 79424 && (row * 584 + col) <= 79640) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 79641 && (row * 584 + col) <= 79887) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 79888 && (row * 584 + col) <= 79930) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 79931 && (row * 584 + col) <= 80007) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 80008 && (row * 584 + col) <= 80224) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 80225 && (row * 584 + col) <= 80472) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 80473 && (row * 584 + col) <= 80513) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 80514 && (row * 584 + col) <= 80591) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 80592 && (row * 584 + col) <= 80808) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 80809 && (row * 584 + col) <= 81057) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 81058 && (row * 584 + col) <= 81096) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 81097 && (row * 584 + col) <= 81175) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 81176 && (row * 584 + col) <= 81392) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 81393 && (row * 584 + col) <= 81642) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 81643 && (row * 584 + col) <= 81679) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 81680 && (row * 584 + col) <= 81759) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 81760 && (row * 584 + col) <= 81976) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 81977 && (row * 584 + col) <= 82228) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 82229 && (row * 584 + col) <= 82261) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 82262 && (row * 584 + col) <= 82343) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 82344 && (row * 584 + col) <= 82560) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 82561 && (row * 584 + col) <= 82814) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 82815 && (row * 584 + col) <= 82843) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 82844 && (row * 584 + col) <= 82927) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 82928 && (row * 584 + col) <= 83144) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 83145 && (row * 584 + col) <= 83400) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 83401 && (row * 584 + col) <= 83425) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 83426 && (row * 584 + col) <= 83511) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 83512 && (row * 584 + col) <= 83728) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 83729 && (row * 584 + col) <= 83987) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 83988 && (row * 584 + col) <= 84006) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 84007 && (row * 584 + col) <= 84095) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 84096 && (row * 584 + col) <= 84312) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 84313 && (row * 584 + col) <= 84575) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 84576 && (row * 584 + col) <= 84586) color_data <= 12'b011111111001; else
        if ((row * 584 + col) >= 84587 && (row * 584 + col) <= 84679) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 84680 && (row * 584 + col) <= 84896) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 84897 && (row * 584 + col) <= 85263) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 85264 && (row * 584 + col) <= 85480) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 85481 && (row * 584 + col) <= 85847) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 85848 && (row * 584 + col) <= 86064) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 86065 && (row * 584 + col) <= 86431) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 86432 && (row * 584 + col) <= 86648) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 86649 && (row * 584 + col) <= 87015) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 87016 && (row * 584 + col) <= 87232) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 87233 && (row * 584 + col) <= 87599) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 87600 && (row * 584 + col) <= 87816) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 87817 && (row * 584 + col) <= 88183) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 88184 && (row * 584 + col) <= 88400) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 88401 && (row * 584 + col) <= 88767) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 88768 && (row * 584 + col) <= 88984) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 88985 && (row * 584 + col) <= 89351) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 89352 && (row * 584 + col) <= 89568) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 89569 && (row * 584 + col) <= 89935) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 89936 && (row * 584 + col) <= 90152) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 90153 && (row * 584 + col) <= 90519) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 90520 && (row * 584 + col) <= 90736) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 90737 && (row * 584 + col) <= 91103) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 91104 && (row * 584 + col) <= 91320) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 91321 && (row * 584 + col) <= 91687) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 91688 && (row * 584 + col) <= 91904) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 91905 && (row * 584 + col) <= 92271) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 92272 && (row * 584 + col) <= 92488) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 92489 && (row * 584 + col) <= 92855) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 92856 && (row * 584 + col) <= 93072) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 93073 && (row * 584 + col) <= 93439) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 93440 && (row * 584 + col) <= 93656) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 93657 && (row * 584 + col) <= 94023) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 94024 && (row * 584 + col) <= 94240) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 94241 && (row * 584 + col) <= 94607) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 94608 && (row * 584 + col) <= 94824) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 94825 && (row * 584 + col) <= 95191) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 95192 && (row * 584 + col) <= 95408) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 95409 && (row * 584 + col) <= 95775) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 95776 && (row * 584 + col) <= 95992) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 95993 && (row * 584 + col) <= 96359) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 96360 && (row * 584 + col) <= 96576) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 96577 && (row * 584 + col) <= 96943) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 96944 && (row * 584 + col) <= 97160) color_data <= 12'b111000010010; else
        if ((row * 584 + col) >= 97161 && (row * 584 + col) < 97528) color_data <= 12'b111111111111; else
        color_data <= 12'b000000000000;
    end
endmodule
