`timescale 1ns / 1ps
module player_rom (
    input wire clk,
    input wire [6:0] row,
    input wire [6:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 100 + col) >= 0 && (row * 100 + col) <= 140) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 141 && (row * 100 + col) <= 155) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 156 && (row * 100 + col) <= 240) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 241 && (row * 100 + col) <= 255) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 256 && (row * 100 + col) <= 333) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 334 && (row * 100 + col) <= 362) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 363 && (row * 100 + col) <= 433) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 434 && (row * 100 + col) <= 462) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 463 && (row * 100 + col) <= 533) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 534 && (row * 100 + col) <= 562) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 563 && (row * 100 + col) <= 631) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 632 && (row * 100 + col) <= 667) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 668 && (row * 100 + col) <= 731) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 732 && (row * 100 + col) <= 767) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 768 && (row * 100 + col) <= 826) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 827 && (row * 100 + col) <= 828) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 829 && (row * 100 + col) <= 867) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 868 && (row * 100 + col) <= 870) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 871 && (row * 100 + col) <= 926) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 927 && (row * 100 + col) <= 928) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 929 && (row * 100 + col) <= 967) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 968 && (row * 100 + col) <= 970) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 971 && (row * 100 + col) <= 1026) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1027 && (row * 100 + col) <= 1028) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1029 && (row * 100 + col) <= 1031) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1032 && (row * 100 + col) <= 1036) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1037 && (row * 100 + col) <= 1043) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1044 && (row * 100 + col) <= 1053) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1054 && (row * 100 + col) <= 1058) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1059 && (row * 100 + col) <= 1065) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1066 && (row * 100 + col) <= 1067) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1068 && (row * 100 + col) <= 1070) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1071 && (row * 100 + col) <= 1126) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1127 && (row * 100 + col) <= 1128) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1129 && (row * 100 + col) <= 1131) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1132 && (row * 100 + col) <= 1136) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1137 && (row * 100 + col) <= 1143) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1144 && (row * 100 + col) <= 1153) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1154 && (row * 100 + col) <= 1158) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1159 && (row * 100 + col) <= 1165) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1166 && (row * 100 + col) <= 1167) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1168 && (row * 100 + col) <= 1170) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1171 && (row * 100 + col) <= 1226) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1227 && (row * 100 + col) <= 1228) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1229 && (row * 100 + col) <= 1231) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1232 && (row * 100 + col) <= 1236) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1237 && (row * 100 + col) <= 1243) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1244 && (row * 100 + col) <= 1253) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1254 && (row * 100 + col) <= 1258) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1259 && (row * 100 + col) <= 1265) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1266 && (row * 100 + col) <= 1267) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1268 && (row * 100 + col) <= 1270) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1271 && (row * 100 + col) <= 1326) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1327 && (row * 100 + col) <= 1331) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1332 && (row * 100 + col) <= 1336) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1337 && (row * 100 + col) <= 1340) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1341 && (row * 100 + col) <= 1343) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1344 && (row * 100 + col) <= 1350) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1351 && (row * 100 + col) <= 1355) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1356 && (row * 100 + col) <= 1358) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1359 && (row * 100 + col) <= 1360) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1361 && (row * 100 + col) <= 1362) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1363 && (row * 100 + col) <= 1365) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1366 && (row * 100 + col) <= 1372) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1373 && (row * 100 + col) <= 1426) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1427 && (row * 100 + col) <= 1431) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1432 && (row * 100 + col) <= 1436) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1437 && (row * 100 + col) <= 1440) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1441 && (row * 100 + col) <= 1443) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1444 && (row * 100 + col) <= 1450) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1451 && (row * 100 + col) <= 1455) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1456 && (row * 100 + col) <= 1458) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1459 && (row * 100 + col) <= 1460) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1461 && (row * 100 + col) <= 1462) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1463 && (row * 100 + col) <= 1465) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1466 && (row * 100 + col) <= 1472) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1473 && (row * 100 + col) <= 1523) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1524 && (row * 100 + col) <= 1533) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1534 && (row * 100 + col) <= 1536) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1537 && (row * 100 + col) <= 1538) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1539 && (row * 100 + col) <= 1540) color_data <= 12'b001101001100; else
        if ((row * 100 + col) >= 1541 && (row * 100 + col) <= 1553) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1554 && (row * 100 + col) <= 1558) color_data <= 12'b001101001100; else
        if ((row * 100 + col) >= 1559 && (row * 100 + col) <= 1562) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1563 && (row * 100 + col) <= 1572) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1573 && (row * 100 + col) <= 1623) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1624 && (row * 100 + col) <= 1633) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1634 && (row * 100 + col) <= 1636) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1637 && (row * 100 + col) <= 1638) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1639 && (row * 100 + col) <= 1640) color_data <= 12'b001101001100; else
        if ((row * 100 + col) >= 1641 && (row * 100 + col) <= 1653) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1654 && (row * 100 + col) <= 1658) color_data <= 12'b001101001100; else
        if ((row * 100 + col) >= 1659 && (row * 100 + col) <= 1662) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1663 && (row * 100 + col) <= 1672) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1673 && (row * 100 + col) <= 1723) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1724 && (row * 100 + col) <= 1736) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1737 && (row * 100 + col) <= 1743) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1744 && (row * 100 + col) <= 1750) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1751 && (row * 100 + col) <= 1753) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1754 && (row * 100 + col) <= 1758) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1759 && (row * 100 + col) <= 1762) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1763 && (row * 100 + col) <= 1772) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1773 && (row * 100 + col) <= 1823) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1824 && (row * 100 + col) <= 1836) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1837 && (row * 100 + col) <= 1843) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1844 && (row * 100 + col) <= 1850) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1851 && (row * 100 + col) <= 1853) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1854 && (row * 100 + col) <= 1858) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1859 && (row * 100 + col) <= 1862) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1863 && (row * 100 + col) <= 1872) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1873 && (row * 100 + col) <= 1923) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 1924 && (row * 100 + col) <= 1936) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1937 && (row * 100 + col) <= 1943) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1944 && (row * 100 + col) <= 1950) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1951 && (row * 100 + col) <= 1953) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1954 && (row * 100 + col) <= 1958) color_data <= 12'b110011001100; else
        if ((row * 100 + col) >= 1959 && (row * 100 + col) <= 1962) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 1963 && (row * 100 + col) <= 1972) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 1973 && (row * 100 + col) <= 2021) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2022 && (row * 100 + col) <= 2053) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2054 && (row * 100 + col) <= 2058) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 2059 && (row * 100 + col) <= 2072) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2073 && (row * 100 + col) <= 2121) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2122 && (row * 100 + col) <= 2153) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2154 && (row * 100 + col) <= 2158) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 2159 && (row * 100 + col) <= 2172) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2173 && (row * 100 + col) <= 2221) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2222 && (row * 100 + col) <= 2272) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2273 && (row * 100 + col) <= 2321) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2322 && (row * 100 + col) <= 2372) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2373 && (row * 100 + col) <= 2421) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2422 && (row * 100 + col) <= 2472) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2473 && (row * 100 + col) <= 2521) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2522 && (row * 100 + col) <= 2572) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2573 && (row * 100 + col) <= 2621) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2622 && (row * 100 + col) <= 2672) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2673 && (row * 100 + col) <= 2723) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2724 && (row * 100 + col) <= 2760) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2761 && (row * 100 + col) <= 2762) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 2763 && (row * 100 + col) <= 2772) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2773 && (row * 100 + col) <= 2823) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2824 && (row * 100 + col) <= 2860) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2861 && (row * 100 + col) <= 2862) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 2863 && (row * 100 + col) <= 2872) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2873 && (row * 100 + col) <= 2923) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 2924 && (row * 100 + col) <= 2933) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2934 && (row * 100 + col) <= 2936) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 2937 && (row * 100 + col) <= 2958) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2959 && (row * 100 + col) <= 2962) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 2963 && (row * 100 + col) <= 2972) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 2973 && (row * 100 + col) <= 3023) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3024 && (row * 100 + col) <= 3033) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3034 && (row * 100 + col) <= 3036) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3037 && (row * 100 + col) <= 3058) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3059 && (row * 100 + col) <= 3062) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3063 && (row * 100 + col) <= 3072) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3073 && (row * 100 + col) <= 3126) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3127 && (row * 100 + col) <= 3133) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3134 && (row * 100 + col) <= 3140) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3141 && (row * 100 + col) <= 3158) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3159 && (row * 100 + col) <= 3160) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3161 && (row * 100 + col) <= 3172) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3173 && (row * 100 + col) <= 3226) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3227 && (row * 100 + col) <= 3233) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3234 && (row * 100 + col) <= 3240) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3241 && (row * 100 + col) <= 3258) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3259 && (row * 100 + col) <= 3260) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3261 && (row * 100 + col) <= 3272) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3273 && (row * 100 + col) <= 3326) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3327 && (row * 100 + col) <= 3333) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3334 && (row * 100 + col) <= 3340) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3341 && (row * 100 + col) <= 3358) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3359 && (row * 100 + col) <= 3360) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3361 && (row * 100 + col) <= 3372) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3373 && (row * 100 + col) <= 3426) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3427 && (row * 100 + col) <= 3438) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3439 && (row * 100 + col) <= 3445) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3446 && (row * 100 + col) <= 3453) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3454 && (row * 100 + col) <= 3458) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3459 && (row * 100 + col) <= 3470) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3471 && (row * 100 + col) <= 3526) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3527 && (row * 100 + col) <= 3538) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3539 && (row * 100 + col) <= 3545) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3546 && (row * 100 + col) <= 3553) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3554 && (row * 100 + col) <= 3558) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3559 && (row * 100 + col) <= 3570) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3571 && (row * 100 + col) <= 3628) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3629 && (row * 100 + col) <= 3640) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3641 && (row * 100 + col) <= 3658) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3659 && (row * 100 + col) <= 3667) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3668 && (row * 100 + col) <= 3728) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3729 && (row * 100 + col) <= 3740) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3741 && (row * 100 + col) <= 3758) color_data <= 12'b000000000000; else
        if ((row * 100 + col) >= 3759 && (row * 100 + col) <= 3767) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3768 && (row * 100 + col) <= 3831) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3832 && (row * 100 + col) <= 3865) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3866 && (row * 100 + col) <= 3931) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 3932 && (row * 100 + col) <= 3965) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 3966 && (row * 100 + col) <= 4031) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4032 && (row * 100 + col) <= 4065) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4066 && (row * 100 + col) <= 4133) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4134 && (row * 100 + col) <= 4162) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4163 && (row * 100 + col) <= 4233) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4234 && (row * 100 + col) <= 4262) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4263 && (row * 100 + col) <= 4340) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4341 && (row * 100 + col) <= 4355) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4356 && (row * 100 + col) <= 4440) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4441 && (row * 100 + col) <= 4455) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4456 && (row * 100 + col) <= 4516) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4517 && (row * 100 + col) <= 4523) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4524 && (row * 100 + col) <= 4540) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4541 && (row * 100 + col) <= 4555) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4556 && (row * 100 + col) <= 4616) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4617 && (row * 100 + col) <= 4623) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4624 && (row * 100 + col) <= 4640) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4641 && (row * 100 + col) <= 4655) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4656 && (row * 100 + col) <= 4716) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4717 && (row * 100 + col) <= 4723) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4724 && (row * 100 + col) <= 4740) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4741 && (row * 100 + col) <= 4755) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4756 && (row * 100 + col) <= 4804) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4805 && (row * 100 + col) <= 4833) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4834 && (row * 100 + col) <= 4838) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4839 && (row * 100 + col) <= 4858) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4859 && (row * 100 + col) <= 4862) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4863 && (row * 100 + col) <= 4892) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4893 && (row * 100 + col) <= 4904) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4905 && (row * 100 + col) <= 4933) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4934 && (row * 100 + col) <= 4938) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4939 && (row * 100 + col) <= 4958) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4959 && (row * 100 + col) <= 4962) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 4963 && (row * 100 + col) <= 4992) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 4993 && (row * 100 + col) <= 5001) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5002 && (row * 100 + col) <= 5094) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5095 && (row * 100 + col) <= 5101) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5102 && (row * 100 + col) <= 5194) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5195 && (row * 100 + col) <= 5201) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5202 && (row * 100 + col) <= 5297) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5298 && (row * 100 + col) <= 5301) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5302 && (row * 100 + col) <= 5397) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5398 && (row * 100 + col) <= 5401) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5402 && (row * 100 + col) <= 5497) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5498 && (row * 100 + col) <= 5501) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5502 && (row * 100 + col) <= 5597) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5598 && (row * 100 + col) <= 5601) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5602 && (row * 100 + col) <= 5697) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5698 && (row * 100 + col) <= 5706) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5707 && (row * 100 + col) <= 5731) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5732 && (row * 100 + col) <= 5736) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5737 && (row * 100 + col) <= 5794) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5795 && (row * 100 + col) <= 5806) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5807 && (row * 100 + col) <= 5831) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5832 && (row * 100 + col) <= 5836) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5837 && (row * 100 + col) <= 5894) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5895 && (row * 100 + col) <= 5933) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5934 && (row * 100 + col) <= 5962) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5963 && (row * 100 + col) <= 5965) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 5966 && (row * 100 + col) <= 5989) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 5990 && (row * 100 + col) <= 6033) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6034 && (row * 100 + col) <= 6062) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6063 && (row * 100 + col) <= 6065) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6066 && (row * 100 + col) <= 6089) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6090 && (row * 100 + col) <= 6133) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6134 && (row * 100 + col) <= 6162) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6163 && (row * 100 + col) <= 6233) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6234 && (row * 100 + col) <= 6262) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6263 && (row * 100 + col) <= 6333) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6334 && (row * 100 + col) <= 6362) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6363 && (row * 100 + col) <= 6436) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6437 && (row * 100 + col) <= 6462) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6463 && (row * 100 + col) <= 6536) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6537 && (row * 100 + col) <= 6562) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6563 && (row * 100 + col) <= 6636) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6637 && (row * 100 + col) <= 6662) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6663 && (row * 100 + col) <= 6736) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6737 && (row * 100 + col) <= 6762) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6763 && (row * 100 + col) <= 6836) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6837 && (row * 100 + col) <= 6860) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6861 && (row * 100 + col) <= 6936) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 6937 && (row * 100 + col) <= 6960) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 6961 && (row * 100 + col) <= 7036) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7037 && (row * 100 + col) <= 7060) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7061 && (row * 100 + col) <= 7136) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7137 && (row * 100 + col) <= 7160) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7161 && (row * 100 + col) <= 7236) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7237 && (row * 100 + col) <= 7260) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7261 && (row * 100 + col) <= 7338) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7339 && (row * 100 + col) <= 7358) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7359 && (row * 100 + col) <= 7438) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7439 && (row * 100 + col) <= 7458) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7459 && (row * 100 + col) <= 7536) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7537 && (row * 100 + col) <= 7560) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7561 && (row * 100 + col) <= 7636) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7637 && (row * 100 + col) <= 7660) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7661 && (row * 100 + col) <= 7736) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7737 && (row * 100 + col) <= 7760) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7761 && (row * 100 + col) <= 7836) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7837 && (row * 100 + col) <= 7843) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7844 && (row * 100 + col) <= 7853) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7854 && (row * 100 + col) <= 7862) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7863 && (row * 100 + col) <= 7936) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7937 && (row * 100 + col) <= 7943) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7944 && (row * 100 + col) <= 7953) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 7954 && (row * 100 + col) <= 7962) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 7963 && (row * 100 + col) <= 8033) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8034 && (row * 100 + col) <= 8045) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8046 && (row * 100 + col) <= 8053) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8054 && (row * 100 + col) <= 8062) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8063 && (row * 100 + col) <= 8133) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8134 && (row * 100 + col) <= 8145) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8146 && (row * 100 + col) <= 8153) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8154 && (row * 100 + col) <= 8162) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8163 && (row * 100 + col) <= 8233) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8234 && (row * 100 + col) <= 8245) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8246 && (row * 100 + col) <= 8253) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8254 && (row * 100 + col) <= 8262) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8263 && (row * 100 + col) <= 8333) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8334 && (row * 100 + col) <= 8345) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8346 && (row * 100 + col) <= 8353) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8354 && (row * 100 + col) <= 8362) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8363 && (row * 100 + col) <= 8433) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8434 && (row * 100 + col) <= 8445) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8446 && (row * 100 + col) <= 8453) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8454 && (row * 100 + col) <= 8462) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8463 && (row * 100 + col) <= 8533) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8534 && (row * 100 + col) <= 8545) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8546 && (row * 100 + col) <= 8553) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8554 && (row * 100 + col) <= 8562) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8563 && (row * 100 + col) <= 8633) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8634 && (row * 100 + col) <= 8645) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8646 && (row * 100 + col) <= 8653) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8654 && (row * 100 + col) <= 8662) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8663 && (row * 100 + col) <= 8733) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8734 && (row * 100 + col) <= 8745) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8746 && (row * 100 + col) <= 8753) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8754 && (row * 100 + col) <= 8762) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8763 && (row * 100 + col) <= 8833) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8834 && (row * 100 + col) <= 8845) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8846 && (row * 100 + col) <= 8853) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8854 && (row * 100 + col) <= 8862) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8863 && (row * 100 + col) <= 8933) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8934 && (row * 100 + col) <= 8945) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8946 && (row * 100 + col) <= 8953) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 8954 && (row * 100 + col) <= 8962) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 8963 && (row * 100 + col) <= 9033) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9034 && (row * 100 + col) <= 9045) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9046 && (row * 100 + col) <= 9053) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9054 && (row * 100 + col) <= 9062) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9063 && (row * 100 + col) <= 9133) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9134 && (row * 100 + col) <= 9145) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9146 && (row * 100 + col) <= 9153) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9154 && (row * 100 + col) <= 9162) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9163 && (row * 100 + col) <= 9236) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9237 && (row * 100 + col) <= 9243) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9244 && (row * 100 + col) <= 9253) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9254 && (row * 100 + col) <= 9262) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9263 && (row * 100 + col) <= 9336) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9337 && (row * 100 + col) <= 9343) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9344 && (row * 100 + col) <= 9353) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9354 && (row * 100 + col) <= 9362) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9363 && (row * 100 + col) <= 9436) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9437 && (row * 100 + col) <= 9443) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9444 && (row * 100 + col) <= 9453) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9454 && (row * 100 + col) <= 9462) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9463 && (row * 100 + col) <= 9536) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9537 && (row * 100 + col) <= 9543) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9544 && (row * 100 + col) <= 9553) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9554 && (row * 100 + col) <= 9562) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9563 && (row * 100 + col) <= 9655) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9656 && (row * 100 + col) <= 9660) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9661 && (row * 100 + col) <= 9755) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9756 && (row * 100 + col) <= 9760) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9761 && (row * 100 + col) <= 9855) color_data <= 12'b111111111111; else
        if ((row * 100 + col) >= 9856 && (row * 100 + col) <= 9860) color_data <= 12'b111011101011; else
        if ((row * 100 + col) >= 9861 && (row * 100 + col) < 10000) color_data <= 12'b111111111111; else
        color_data <= 12'b000000000000;
    end
endmodule
