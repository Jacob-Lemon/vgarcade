module three_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "distributed" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		10'b0000100101: color_data = 12'b000000000000;
		10'b0000100110: color_data = 12'b000000000000;
		10'b0000100111: color_data = 12'b000000000000;
		10'b0000101000: color_data = 12'b000000000000;
		10'b0000101001: color_data = 12'b000000000000;
		10'b0000101010: color_data = 12'b000000000000;
		10'b0000101011: color_data = 12'b000000000000;
		10'b0000101100: color_data = 12'b000000000000;
		10'b0000101101: color_data = 12'b000000000000;
		10'b0000101110: color_data = 12'b000000000000;
		10'b0000101111: color_data = 12'b000000000000;
		10'b0000110000: color_data = 12'b000000000000;
		10'b0001000010: color_data = 12'b000000000000;
		10'b0001000011: color_data = 12'b000000000000;
		10'b0001000100: color_data = 12'b000000000000;
		10'b0001000101: color_data = 12'b000000000000;
		10'b0001000110: color_data = 12'b000000000000;
		10'b0001000111: color_data = 12'b000000000000;
		10'b0001001000: color_data = 12'b000000000000;
		10'b0001001001: color_data = 12'b000000000000;
		10'b0001001010: color_data = 12'b000000000000;
		10'b0001001011: color_data = 12'b000000000000;
		10'b0001001100: color_data = 12'b000000000000;
		10'b0001001101: color_data = 12'b000000000000;
		10'b0001001110: color_data = 12'b000000000000;
		10'b0001001111: color_data = 12'b000000000000;
		10'b0001010000: color_data = 12'b000000000000;
		10'b0001010001: color_data = 12'b000000000000;
		10'b0001010010: color_data = 12'b000000000000;
		10'b0001100001: color_data = 12'b000000000000;
		10'b0001100010: color_data = 12'b000000000000;
		10'b0001100011: color_data = 12'b000000000000;
		10'b0001100100: color_data = 12'b000000000000;
		10'b0001100101: color_data = 12'b000000000000;
		10'b0001100110: color_data = 12'b000000000000;
		10'b0001100111: color_data = 12'b000000000000;
		10'b0001101000: color_data = 12'b000000000000;
		10'b0001101001: color_data = 12'b000000000000;
		10'b0001101010: color_data = 12'b000000000000;
		10'b0001101011: color_data = 12'b000000000000;
		10'b0001101100: color_data = 12'b000000000000;
		10'b0001101101: color_data = 12'b000000000000;
		10'b0001101110: color_data = 12'b000000000000;
		10'b0001101111: color_data = 12'b000000000000;
		10'b0001110000: color_data = 12'b000000000000;
		10'b0001110001: color_data = 12'b000000000000;
		10'b0001110010: color_data = 12'b000000000000;
		10'b0001110011: color_data = 12'b000000000000;
		10'b0010000001: color_data = 12'b000000000000;
		10'b0010000010: color_data = 12'b000000000000;
		10'b0010000011: color_data = 12'b000000000000;
		10'b0010000100: color_data = 12'b000000000000;
		10'b0010000101: color_data = 12'b000000000000;
		10'b0010000110: color_data = 12'b000000000000;
		10'b0010000111: color_data = 12'b000000000000;
		10'b0010001110: color_data = 12'b000000000000;
		10'b0010001111: color_data = 12'b000000000000;
		10'b0010010000: color_data = 12'b000000000000;
		10'b0010010001: color_data = 12'b000000000000;
		10'b0010010010: color_data = 12'b000000000000;
		10'b0010010011: color_data = 12'b000000000000;
		10'b0010010100: color_data = 12'b000000000000;
		10'b0010100001: color_data = 12'b000000000000;
		10'b0010100010: color_data = 12'b000000000000;
		10'b0010100011: color_data = 12'b000000000000;
		10'b0010100100: color_data = 12'b000000000000;
		10'b0010110000: color_data = 12'b000000000000;
		10'b0010110001: color_data = 12'b000000000000;
		10'b0010110010: color_data = 12'b000000000000;
		10'b0010110011: color_data = 12'b000000000000;
		10'b0010110100: color_data = 12'b000000000000;
		10'b0010110101: color_data = 12'b000000000000;
		10'b0011010001: color_data = 12'b000000000000;
		10'b0011010010: color_data = 12'b000000000000;
		10'b0011010011: color_data = 12'b000000000000;
		10'b0011010100: color_data = 12'b000000000000;
		10'b0011010101: color_data = 12'b000000000000;
		10'b0011110010: color_data = 12'b000000000000;
		10'b0011110011: color_data = 12'b000000000000;
		10'b0011110100: color_data = 12'b000000000000;
		10'b0011110101: color_data = 12'b000000000000;
		10'b0011110110: color_data = 12'b000000000000;
		10'b0100010011: color_data = 12'b000000000000;
		10'b0100010100: color_data = 12'b000000000000;
		10'b0100010101: color_data = 12'b000000000000;
		10'b0100010110: color_data = 12'b000000000000;
		10'b0100110011: color_data = 12'b000000000000;
		10'b0100110100: color_data = 12'b000000000000;
		10'b0100110101: color_data = 12'b000000000000;
		10'b0100110110: color_data = 12'b000000000000;
		10'b0100110111: color_data = 12'b000000000000;
		10'b0101010011: color_data = 12'b000000000000;
		10'b0101010100: color_data = 12'b000000000000;
		10'b0101010101: color_data = 12'b000000000000;
		10'b0101010110: color_data = 12'b000000000000;
		10'b0101010111: color_data = 12'b000000000000;
		10'b0101110011: color_data = 12'b000000000000;
		10'b0101110100: color_data = 12'b000000000000;
		10'b0101110101: color_data = 12'b000000000000;
		10'b0101110110: color_data = 12'b000000000000;
		10'b0101110111: color_data = 12'b000000000000;
		10'b0110001111: color_data = 12'b000000000000;
		10'b0110010000: color_data = 12'b000000000000;
		10'b0110010001: color_data = 12'b000000000000;
		10'b0110010010: color_data = 12'b000000000000;
		10'b0110010011: color_data = 12'b000000000000;
		10'b0110010100: color_data = 12'b000000000000;
		10'b0110010101: color_data = 12'b000000000000;
		10'b0110010110: color_data = 12'b000000000000;
		10'b0110101011: color_data = 12'b000000000000;
		10'b0110101100: color_data = 12'b000000000000;
		10'b0110101101: color_data = 12'b000000000000;
		10'b0110101110: color_data = 12'b000000000000;
		10'b0110101111: color_data = 12'b000000000000;
		10'b0110110000: color_data = 12'b000000000000;
		10'b0110110001: color_data = 12'b000000000000;
		10'b0110110010: color_data = 12'b000000000000;
		10'b0110110011: color_data = 12'b000000000000;
		10'b0110110100: color_data = 12'b000000000000;
		10'b0110110101: color_data = 12'b000000000000;
		10'b0111001011: color_data = 12'b000000000000;
		10'b0111001100: color_data = 12'b000000000000;
		10'b0111001101: color_data = 12'b000000000000;
		10'b0111001110: color_data = 12'b000000000000;
		10'b0111001111: color_data = 12'b000000000000;
		10'b0111010000: color_data = 12'b000000000000;
		10'b0111010001: color_data = 12'b000000000000;
		10'b0111010010: color_data = 12'b000000000000;
		10'b0111010011: color_data = 12'b000000000000;
		10'b0111010100: color_data = 12'b000000000000;
		10'b0111010101: color_data = 12'b000000000000;
		10'b0111101011: color_data = 12'b000000000000;
		10'b0111101100: color_data = 12'b000000000000;
		10'b0111101101: color_data = 12'b000000000000;
		10'b0111101110: color_data = 12'b000000000000;
		10'b0111101111: color_data = 12'b000000000000;
		10'b0111110000: color_data = 12'b000000000000;
		10'b0111110001: color_data = 12'b000000000000;
		10'b0111110010: color_data = 12'b000000000000;
		10'b0111110011: color_data = 12'b000000000000;
		10'b0111110100: color_data = 12'b000000000000;
		10'b0111110101: color_data = 12'b000000000000;
		10'b0111110110: color_data = 12'b000000000000;
		10'b1000001011: color_data = 12'b000000000000;
		10'b1000001100: color_data = 12'b000000000000;
		10'b1000001101: color_data = 12'b000000000000;
		10'b1000001110: color_data = 12'b000000000000;
		10'b1000001111: color_data = 12'b000000000000;
		10'b1000010000: color_data = 12'b000000000000;
		10'b1000010001: color_data = 12'b000000000000;
		10'b1000010010: color_data = 12'b000000000000;
		10'b1000010011: color_data = 12'b000000000000;
		10'b1000010100: color_data = 12'b000000000000;
		10'b1000010101: color_data = 12'b000000000000;
		10'b1000010110: color_data = 12'b000000000000;
		10'b1000110011: color_data = 12'b000000000000;
		10'b1000110100: color_data = 12'b000000000000;
		10'b1000110101: color_data = 12'b000000000000;
		10'b1000110110: color_data = 12'b000000000000;
		10'b1001010100: color_data = 12'b000000000000;
		10'b1001010101: color_data = 12'b000000000000;
		10'b1001010110: color_data = 12'b000000000000;
		10'b1001010111: color_data = 12'b000000000000;
		10'b1001110100: color_data = 12'b000000000000;
		10'b1001110101: color_data = 12'b000000000000;
		10'b1001110110: color_data = 12'b000000000000;
		10'b1001110111: color_data = 12'b000000000000;
		10'b1010010100: color_data = 12'b000000000000;
		10'b1010010101: color_data = 12'b000000000000;
		10'b1010010110: color_data = 12'b000000000000;
		10'b1010010111: color_data = 12'b000000000000;
		10'b1010110011: color_data = 12'b000000000000;
		10'b1010110100: color_data = 12'b000000000000;
		10'b1010110101: color_data = 12'b000000000000;
		10'b1010110110: color_data = 12'b000000000000;
		10'b1010110111: color_data = 12'b000000000000;
		10'b1011010011: color_data = 12'b000000000000;
		10'b1011010100: color_data = 12'b000000000000;
		10'b1011010101: color_data = 12'b000000000000;
		10'b1011010110: color_data = 12'b000000000000;
		10'b1011110010: color_data = 12'b000000000000;
		10'b1011110011: color_data = 12'b000000000000;
		10'b1011110100: color_data = 12'b000000000000;
		10'b1011110101: color_data = 12'b000000000000;
		10'b1011110110: color_data = 12'b000000000000;
		10'b1100000010: color_data = 12'b000000000000;
		10'b1100000011: color_data = 12'b000000000000;
		10'b1100010000: color_data = 12'b000000000000;
		10'b1100010001: color_data = 12'b000000000000;
		10'b1100010010: color_data = 12'b000000000000;
		10'b1100010011: color_data = 12'b000000000000;
		10'b1100010100: color_data = 12'b000000000000;
		10'b1100010101: color_data = 12'b000000000000;
		10'b1100100010: color_data = 12'b000000000000;
		10'b1100100011: color_data = 12'b000000000000;
		10'b1100100100: color_data = 12'b000000000000;
		10'b1100101100: color_data = 12'b000000000000;
		10'b1100101101: color_data = 12'b000000000000;
		10'b1100101110: color_data = 12'b000000000000;
		10'b1100101111: color_data = 12'b000000000000;
		10'b1100110000: color_data = 12'b000000000000;
		10'b1100110001: color_data = 12'b000000000000;
		10'b1100110010: color_data = 12'b000000000000;
		10'b1100110011: color_data = 12'b000000000000;
		10'b1100110100: color_data = 12'b000000000000;
		10'b1100110101: color_data = 12'b000000000000;
		10'b1101000010: color_data = 12'b000000000000;
		10'b1101000011: color_data = 12'b000000000000;
		10'b1101000100: color_data = 12'b000000000000;
		10'b1101000101: color_data = 12'b000000000000;
		10'b1101000110: color_data = 12'b000000000000;
		10'b1101000111: color_data = 12'b000000000000;
		10'b1101001000: color_data = 12'b000000000000;
		10'b1101001001: color_data = 12'b000000000000;
		10'b1101001010: color_data = 12'b000000000000;
		10'b1101001011: color_data = 12'b000000000000;
		10'b1101001100: color_data = 12'b000000000000;
		10'b1101001101: color_data = 12'b000000000000;
		10'b1101001110: color_data = 12'b000000000000;
		10'b1101001111: color_data = 12'b000000000000;
		10'b1101010000: color_data = 12'b000000000000;
		10'b1101010001: color_data = 12'b000000000000;
		10'b1101010010: color_data = 12'b000000000000;
		10'b1101010011: color_data = 12'b000000000000;
		10'b1101010100: color_data = 12'b000000000000;
		10'b1101100010: color_data = 12'b000000000000;
		10'b1101100011: color_data = 12'b000000000000;
		10'b1101100100: color_data = 12'b000000000000;
		10'b1101100101: color_data = 12'b000000000000;
		10'b1101100110: color_data = 12'b000000000000;
		10'b1101100111: color_data = 12'b000000000000;
		10'b1101101000: color_data = 12'b000000000000;
		10'b1101101001: color_data = 12'b000000000000;
		10'b1101101010: color_data = 12'b000000000000;
		10'b1101101011: color_data = 12'b000000000000;
		10'b1101101100: color_data = 12'b000000000000;
		10'b1101101101: color_data = 12'b000000000000;
		10'b1101101110: color_data = 12'b000000000000;
		10'b1101101111: color_data = 12'b000000000000;
		10'b1101110000: color_data = 12'b000000000000;
		10'b1101110001: color_data = 12'b000000000000;
		10'b1101110010: color_data = 12'b000000000000;
		10'b1110000011: color_data = 12'b000000000000;
		10'b1110000100: color_data = 12'b000000000000;
		10'b1110000101: color_data = 12'b000000000000;
		10'b1110000110: color_data = 12'b000000000000;
		10'b1110000111: color_data = 12'b000000000000;
		10'b1110001000: color_data = 12'b000000000000;
		10'b1110001001: color_data = 12'b000000000000;
		10'b1110001010: color_data = 12'b000000000000;
		10'b1110001011: color_data = 12'b000000000000;
		10'b1110001100: color_data = 12'b000000000000;
		10'b1110001101: color_data = 12'b000000000000;
		10'b1110001110: color_data = 12'b000000000000;
        default: color_data = 12'b111111111111;
	endcase
endmodule