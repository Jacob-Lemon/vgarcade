module start_screen_rom (
    input wire clk,
    input wire [8:0] row,
    input wire [9:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 640 + col) >= 0 && (row * 640 + col) <= 12841) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 12842 && (row * 640 + col) <= 12850) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 12851 && (row * 640 + col) <= 13480) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 13481 && (row * 640 + col) <= 13482) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 13483 && (row * 640 + col) <= 13489) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 13490 && (row * 640 + col) <= 13492) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 13493 && (row * 640 + col) <= 14038) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 14039 && (row * 640 + col) <= 14047) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14048 && (row * 640 + col) <= 14115) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 14116 && (row * 640 + col) <= 14117) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 14118 && (row * 640 + col) <= 14119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 14120 && (row * 640 + col) <= 14121) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 14122 && (row * 640 + col) <= 14131) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 14132 && (row * 640 + col) <= 14133) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 14134 && (row * 640 + col) <= 14677) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 14678 && (row * 640 + col) <= 14679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14680 && (row * 640 + col) <= 14686) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 14687 && (row * 640 + col) <= 14689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14690 && (row * 640 + col) <= 14755) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 14756 && (row * 640 + col) <= 14756) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 14757 && (row * 640 + col) <= 14759) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14760 && (row * 640 + col) <= 14760) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 14761 && (row * 640 + col) <= 14766) color_data <= 12'b000110000011; else
        if ((row * 640 + col) >= 14767 && (row * 640 + col) <= 14768) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 14769 && (row * 640 + col) <= 14772) color_data <= 12'b000110000011; else
        if ((row * 640 + col) >= 14773 && (row * 640 + col) <= 14773) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 14774 && (row * 640 + col) <= 14774) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 14775 && (row * 640 + col) <= 15312) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 15313 && (row * 640 + col) <= 15314) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15315 && (row * 640 + col) <= 15316) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 15317 && (row * 640 + col) <= 15318) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15319 && (row * 640 + col) <= 15328) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 15329 && (row * 640 + col) <= 15330) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15331 && (row * 640 + col) <= 15396) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 15397 && (row * 640 + col) <= 15397) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 15398 && (row * 640 + col) <= 15398) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 15399 && (row * 640 + col) <= 15399) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15400 && (row * 640 + col) <= 15401) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 15402 && (row * 640 + col) <= 15413) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 15414 && (row * 640 + col) <= 15415) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15416 && (row * 640 + col) <= 15952) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 15953 && (row * 640 + col) <= 15953) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15954 && (row * 640 + col) <= 15956) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 15957 && (row * 640 + col) <= 15957) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15958 && (row * 640 + col) <= 15963) color_data <= 12'b000110000011; else
        if ((row * 640 + col) >= 15964 && (row * 640 + col) <= 15965) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 15966 && (row * 640 + col) <= 15969) color_data <= 12'b000110000011; else
        if ((row * 640 + col) >= 15970 && (row * 640 + col) <= 15970) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 15971 && (row * 640 + col) <= 15971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 15972 && (row * 640 + col) <= 16036) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 16037 && (row * 640 + col) <= 16037) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16038 && (row * 640 + col) <= 16041) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 16042 && (row * 640 + col) <= 16054) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 16055 && (row * 640 + col) <= 16055) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 16056 && (row * 640 + col) <= 16593) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 16594 && (row * 640 + col) <= 16594) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16595 && (row * 640 + col) <= 16595) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 16596 && (row * 640 + col) <= 16596) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 16597 && (row * 640 + col) <= 16598) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 16599 && (row * 640 + col) <= 16610) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 16611 && (row * 640 + col) <= 16612) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 16613 && (row * 640 + col) <= 16668) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 16669 && (row * 640 + col) <= 16674) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 16675 && (row * 640 + col) <= 16675) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16676 && (row * 640 + col) <= 16676) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 16677 && (row * 640 + col) <= 16677) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16678 && (row * 640 + col) <= 16678) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 16679 && (row * 640 + col) <= 16681) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 16682 && (row * 640 + col) <= 16687) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 16688 && (row * 640 + col) <= 16692) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 16693 && (row * 640 + col) <= 16693) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 16694 && (row * 640 + col) <= 16695) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 16696 && (row * 640 + col) <= 17233) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 17234 && (row * 640 + col) <= 17234) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17235 && (row * 640 + col) <= 17238) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 17239 && (row * 640 + col) <= 17251) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 17252 && (row * 640 + col) <= 17252) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17253 && (row * 640 + col) <= 17306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 17307 && (row * 640 + col) <= 17308) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17309 && (row * 640 + col) <= 17309) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17310 && (row * 640 + col) <= 17314) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 17315 && (row * 640 + col) <= 17316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17317 && (row * 640 + col) <= 17317) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17318 && (row * 640 + col) <= 17318) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17319 && (row * 640 + col) <= 17320) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 17321 && (row * 640 + col) <= 17321) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17322 && (row * 640 + col) <= 17322) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17323 && (row * 640 + col) <= 17326) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 17327 && (row * 640 + col) <= 17332) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17333 && (row * 640 + col) <= 17333) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17334 && (row * 640 + col) <= 17865) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 17866 && (row * 640 + col) <= 17871) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17872 && (row * 640 + col) <= 17874) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17875 && (row * 640 + col) <= 17878) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 17879 && (row * 640 + col) <= 17884) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17885 && (row * 640 + col) <= 17889) color_data <= 12'b000110010100; else
        if ((row * 640 + col) >= 17890 && (row * 640 + col) <= 17890) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17891 && (row * 640 + col) <= 17892) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17893 && (row * 640 + col) <= 17945) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 17946 && (row * 640 + col) <= 17947) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17948 && (row * 640 + col) <= 17955) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 17956 && (row * 640 + col) <= 17957) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17958 && (row * 640 + col) <= 17958) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17959 && (row * 640 + col) <= 17960) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 17961 && (row * 640 + col) <= 17961) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17962 && (row * 640 + col) <= 17967) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 17968 && (row * 640 + col) <= 17968) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 17969 && (row * 640 + col) <= 17969) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 17970 && (row * 640 + col) <= 18503) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 18504 && (row * 640 + col) <= 18505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18506 && (row * 640 + col) <= 18506) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 18507 && (row * 640 + col) <= 18513) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 18514 && (row * 640 + col) <= 18514) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18515 && (row * 640 + col) <= 18515) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 18516 && (row * 640 + col) <= 18517) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 18518 && (row * 640 + col) <= 18518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18519 && (row * 640 + col) <= 18519) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 18520 && (row * 640 + col) <= 18523) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 18524 && (row * 640 + col) <= 18529) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 18530 && (row * 640 + col) <= 18530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18531 && (row * 640 + col) <= 18584) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 18585 && (row * 640 + col) <= 18586) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18587 && (row * 640 + col) <= 18589) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 18590 && (row * 640 + col) <= 18592) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 18593 && (row * 640 + col) <= 18597) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 18598 && (row * 640 + col) <= 18598) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 18599 && (row * 640 + col) <= 18600) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 18601 && (row * 640 + col) <= 18601) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 18602 && (row * 640 + col) <= 18608) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 18609 && (row * 640 + col) <= 18610) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 18611 && (row * 640 + col) <= 18611) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 18612 && (row * 640 + col) <= 19142) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 19143 && (row * 640 + col) <= 19144) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19145 && (row * 640 + col) <= 19154) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 19155 && (row * 640 + col) <= 19155) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 19156 && (row * 640 + col) <= 19157) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 19158 && (row * 640 + col) <= 19158) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 19159 && (row * 640 + col) <= 19164) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 19165 && (row * 640 + col) <= 19165) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19166 && (row * 640 + col) <= 19166) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 19167 && (row * 640 + col) <= 19223) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 19224 && (row * 640 + col) <= 19225) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19226 && (row * 640 + col) <= 19234) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 19235 && (row * 640 + col) <= 19238) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 19239 && (row * 640 + col) <= 19240) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 19241 && (row * 640 + col) <= 19250) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 19251 && (row * 640 + col) <= 19251) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 19252 && (row * 640 + col) <= 19252) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19253 && (row * 640 + col) <= 19781) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 19782 && (row * 640 + col) <= 19783) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19784 && (row * 640 + col) <= 19789) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 19790 && (row * 640 + col) <= 19795) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 19796 && (row * 640 + col) <= 19797) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 19798 && (row * 640 + col) <= 19805) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 19806 && (row * 640 + col) <= 19807) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 19808 && (row * 640 + col) <= 19808) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19809 && (row * 640 + col) <= 19862) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 19863 && (row * 640 + col) <= 19863) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 19864 && (row * 640 + col) <= 19864) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 19865 && (row * 640 + col) <= 19875) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 19876 && (row * 640 + col) <= 19878) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 19879 && (row * 640 + col) <= 19880) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 19881 && (row * 640 + col) <= 19891) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 19892 && (row * 640 + col) <= 19893) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 19894 && (row * 640 + col) <= 20420) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 20421 && (row * 640 + col) <= 20422) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20423 && (row * 640 + col) <= 20431) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 20432 && (row * 640 + col) <= 20435) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 20436 && (row * 640 + col) <= 20437) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 20438 && (row * 640 + col) <= 20447) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 20448 && (row * 640 + col) <= 20448) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 20449 && (row * 640 + col) <= 20449) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20450 && (row * 640 + col) <= 20501) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 20502 && (row * 640 + col) <= 20503) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20504 && (row * 640 + col) <= 20516) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 20517 && (row * 640 + col) <= 20532) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 20533 && (row * 640 + col) <= 20533) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 20534 && (row * 640 + col) <= 20534) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 20535 && (row * 640 + col) <= 21059) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 21060 && (row * 640 + col) <= 21060) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21061 && (row * 640 + col) <= 21061) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 21062 && (row * 640 + col) <= 21072) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 21073 && (row * 640 + col) <= 21075) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 21076 && (row * 640 + col) <= 21077) color_data <= 12'b011101000011; else
        if ((row * 640 + col) >= 21078 && (row * 640 + col) <= 21088) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 21089 && (row * 640 + col) <= 21090) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 21091 && (row * 640 + col) <= 21141) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 21142 && (row * 640 + col) <= 21142) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 21143 && (row * 640 + col) <= 21147) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 21148 && (row * 640 + col) <= 21150) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 21151 && (row * 640 + col) <= 21162) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 21163 && (row * 640 + col) <= 21173) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 21174 && (row * 640 + col) <= 21174) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 21175 && (row * 640 + col) <= 21175) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21176 && (row * 640 + col) <= 21698) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 21699 && (row * 640 + col) <= 21700) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21701 && (row * 640 + col) <= 21713) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 21714 && (row * 640 + col) <= 21729) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 21730 && (row * 640 + col) <= 21730) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 21731 && (row * 640 + col) <= 21731) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21732 && (row * 640 + col) <= 21780) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 21781 && (row * 640 + col) <= 21781) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 21782 && (row * 640 + col) <= 21782) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 21783 && (row * 640 + col) <= 21786) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 21787 && (row * 640 + col) <= 21790) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 21791 && (row * 640 + col) <= 21804) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 21805 && (row * 640 + col) <= 21814) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 21815 && (row * 640 + col) <= 21815) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 21816 && (row * 640 + col) <= 22338) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 22339 && (row * 640 + col) <= 22339) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 22340 && (row * 640 + col) <= 22344) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 22345 && (row * 640 + col) <= 22347) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 22348 && (row * 640 + col) <= 22359) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 22360 && (row * 640 + col) <= 22370) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 22371 && (row * 640 + col) <= 22371) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 22372 && (row * 640 + col) <= 22420) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 22421 && (row * 640 + col) <= 22421) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22422 && (row * 640 + col) <= 22425) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 22426 && (row * 640 + col) <= 22429) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 22430 && (row * 640 + col) <= 22444) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 22445 && (row * 640 + col) <= 22454) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 22455 && (row * 640 + col) <= 22455) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 22456 && (row * 640 + col) <= 22456) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22457 && (row * 640 + col) <= 22977) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 22978 && (row * 640 + col) <= 22978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 22979 && (row * 640 + col) <= 22979) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 22980 && (row * 640 + col) <= 22983) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 22984 && (row * 640 + col) <= 22987) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 22988 && (row * 640 + col) <= 23001) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 23002 && (row * 640 + col) <= 23010) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 23011 && (row * 640 + col) <= 23011) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23012 && (row * 640 + col) <= 23012) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 23013 && (row * 640 + col) <= 23060) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 23061 && (row * 640 + col) <= 23061) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23062 && (row * 640 + col) <= 23065) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 23066 && (row * 640 + col) <= 23068) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 23069 && (row * 640 + col) <= 23085) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 23086 && (row * 640 + col) <= 23095) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 23096 && (row * 640 + col) <= 23096) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23097 && (row * 640 + col) <= 23617) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 23618 && (row * 640 + col) <= 23618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23619 && (row * 640 + col) <= 23622) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 23623 && (row * 640 + col) <= 23626) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 23627 && (row * 640 + col) <= 23641) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 23642 && (row * 640 + col) <= 23651) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 23652 && (row * 640 + col) <= 23652) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 23653 && (row * 640 + col) <= 23700) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 23701 && (row * 640 + col) <= 23701) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23702 && (row * 640 + col) <= 23705) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 23706 && (row * 640 + col) <= 23707) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 23708 && (row * 640 + col) <= 23726) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 23727 && (row * 640 + col) <= 23735) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 23736 && (row * 640 + col) <= 23736) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 23737 && (row * 640 + col) <= 24257) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 24258 && (row * 640 + col) <= 24258) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24259 && (row * 640 + col) <= 24262) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 24263 && (row * 640 + col) <= 24265) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 24266 && (row * 640 + col) <= 24282) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 24283 && (row * 640 + col) <= 24291) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 24292 && (row * 640 + col) <= 24293) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24294 && (row * 640 + col) <= 24340) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 24341 && (row * 640 + col) <= 24341) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24342 && (row * 640 + col) <= 24366) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 24367 && (row * 640 + col) <= 24375) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 24376 && (row * 640 + col) <= 24376) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24377 && (row * 640 + col) <= 24897) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 24898 && (row * 640 + col) <= 24898) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24899 && (row * 640 + col) <= 24902) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 24903 && (row * 640 + col) <= 24904) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 24905 && (row * 640 + col) <= 24923) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 24924 && (row * 640 + col) <= 24932) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 24933 && (row * 640 + col) <= 24933) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24934 && (row * 640 + col) <= 24980) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 24981 && (row * 640 + col) <= 24981) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 24982 && (row * 640 + col) <= 25006) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 25007 && (row * 640 + col) <= 25015) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 25016 && (row * 640 + col) <= 25016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25017 && (row * 640 + col) <= 25537) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 25538 && (row * 640 + col) <= 25538) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25539 && (row * 640 + col) <= 25563) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 25564 && (row * 640 + col) <= 25572) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 25573 && (row * 640 + col) <= 25573) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25574 && (row * 640 + col) <= 25620) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 25621 && (row * 640 + col) <= 25621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25622 && (row * 640 + col) <= 25646) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 25647 && (row * 640 + col) <= 25655) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 25656 && (row * 640 + col) <= 25656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 25657 && (row * 640 + col) <= 26177) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 26178 && (row * 640 + col) <= 26178) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26179 && (row * 640 + col) <= 26203) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 26204 && (row * 640 + col) <= 26212) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 26213 && (row * 640 + col) <= 26213) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26214 && (row * 640 + col) <= 26260) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 26261 && (row * 640 + col) <= 26261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26262 && (row * 640 + col) <= 26262) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 26263 && (row * 640 + col) <= 26286) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 26287 && (row * 640 + col) <= 26295) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 26296 && (row * 640 + col) <= 26296) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26297 && (row * 640 + col) <= 26817) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 26818 && (row * 640 + col) <= 26818) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26819 && (row * 640 + col) <= 26843) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 26844 && (row * 640 + col) <= 26852) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 26853 && (row * 640 + col) <= 26853) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26854 && (row * 640 + col) <= 26901) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 26902 && (row * 640 + col) <= 26902) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 26903 && (row * 640 + col) <= 26926) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 26927 && (row * 640 + col) <= 26935) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 26936 && (row * 640 + col) <= 26936) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 26937 && (row * 640 + col) <= 27457) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 27458 && (row * 640 + col) <= 27458) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27459 && (row * 640 + col) <= 27483) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 27484 && (row * 640 + col) <= 27492) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 27493 && (row * 640 + col) <= 27493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27494 && (row * 640 + col) <= 27541) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 27542 && (row * 640 + col) <= 27543) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 27544 && (row * 640 + col) <= 27566) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 27567 && (row * 640 + col) <= 27575) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 27576 && (row * 640 + col) <= 27576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 27577 && (row * 640 + col) <= 28097) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 28098 && (row * 640 + col) <= 28098) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28099 && (row * 640 + col) <= 28099) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 28100 && (row * 640 + col) <= 28123) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 28124 && (row * 640 + col) <= 28132) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 28133 && (row * 640 + col) <= 28133) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28134 && (row * 640 + col) <= 28182) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 28183 && (row * 640 + col) <= 28183) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28184 && (row * 640 + col) <= 28184) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 28185 && (row * 640 + col) <= 28206) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 28207 && (row * 640 + col) <= 28214) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 28215 && (row * 640 + col) <= 28216) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28217 && (row * 640 + col) <= 28738) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 28739 && (row * 640 + col) <= 28739) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 28740 && (row * 640 + col) <= 28740) color_data <= 12'b110001100001; else
        if ((row * 640 + col) >= 28741 && (row * 640 + col) <= 28763) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 28764 && (row * 640 + col) <= 28772) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 28773 && (row * 640 + col) <= 28773) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28774 && (row * 640 + col) <= 28822) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 28823 && (row * 640 + col) <= 28823) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28824 && (row * 640 + col) <= 28824) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 28825 && (row * 640 + col) <= 28825) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 28826 && (row * 640 + col) <= 28846) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 28847 && (row * 640 + col) <= 28854) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 28855 && (row * 640 + col) <= 28855) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 28856 && (row * 640 + col) <= 29378) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 29379 && (row * 640 + col) <= 29380) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29381 && (row * 640 + col) <= 29403) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 29404 && (row * 640 + col) <= 29411) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 29412 && (row * 640 + col) <= 29413) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29414 && (row * 640 + col) <= 29463) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 29464 && (row * 640 + col) <= 29464) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 29465 && (row * 640 + col) <= 29466) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 29467 && (row * 640 + col) <= 29485) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 29486 && (row * 640 + col) <= 29493) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 29494 && (row * 640 + col) <= 29495) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 29496 && (row * 640 + col) <= 30019) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 30020 && (row * 640 + col) <= 30020) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30021 && (row * 640 + col) <= 30021) color_data <= 12'b110001100001; else
        if ((row * 640 + col) >= 30022 && (row * 640 + col) <= 30043) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 30044 && (row * 640 + col) <= 30051) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 30052 && (row * 640 + col) <= 30052) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30053 && (row * 640 + col) <= 30103) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 30104 && (row * 640 + col) <= 30105) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 30106 && (row * 640 + col) <= 30106) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 30107 && (row * 640 + col) <= 30124) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 30125 && (row * 640 + col) <= 30132) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 30133 && (row * 640 + col) <= 30133) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 30134 && (row * 640 + col) <= 30134) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30135 && (row * 640 + col) <= 30659) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 30660 && (row * 640 + col) <= 30660) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30661 && (row * 640 + col) <= 30661) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 30662 && (row * 640 + col) <= 30662) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 30663 && (row * 640 + col) <= 30682) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 30683 && (row * 640 + col) <= 30690) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 30691 && (row * 640 + col) <= 30692) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30693 && (row * 640 + col) <= 30744) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 30745 && (row * 640 + col) <= 30745) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 30746 && (row * 640 + col) <= 30746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 30747 && (row * 640 + col) <= 30747) color_data <= 12'b101000000000; else
        if ((row * 640 + col) >= 30748 && (row * 640 + col) <= 30763) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 30764 && (row * 640 + col) <= 30771) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 30772 && (row * 640 + col) <= 30773) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 30774 && (row * 640 + col) <= 31300) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 31301 && (row * 640 + col) <= 31301) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 31302 && (row * 640 + col) <= 31303) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 31304 && (row * 640 + col) <= 31321) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 31322 && (row * 640 + col) <= 31330) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 31331 && (row * 640 + col) <= 31331) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31332 && (row * 640 + col) <= 31385) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 31386 && (row * 640 + col) <= 31386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31387 && (row * 640 + col) <= 31387) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 31388 && (row * 640 + col) <= 31389) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 31390 && (row * 640 + col) <= 31402) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 31403 && (row * 640 + col) <= 31410) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 31411 && (row * 640 + col) <= 31412) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31413 && (row * 640 + col) <= 31940) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 31941 && (row * 640 + col) <= 31941) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31942 && (row * 640 + col) <= 31942) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 31943 && (row * 640 + col) <= 31944) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 31945 && (row * 640 + col) <= 31960) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 31961 && (row * 640 + col) <= 31969) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 31970 && (row * 640 + col) <= 31970) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 31971 && (row * 640 + col) <= 31971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 31972 && (row * 640 + col) <= 32026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 32027 && (row * 640 + col) <= 32028) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 32029 && (row * 640 + col) <= 32030) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 32031 && (row * 640 + col) <= 32040) color_data <= 12'b111100000000; else
        if ((row * 640 + col) >= 32041 && (row * 640 + col) <= 32049) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 32050 && (row * 640 + col) <= 32050) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 32051 && (row * 640 + col) <= 32051) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32052 && (row * 640 + col) <= 32581) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 32582 && (row * 640 + col) <= 32583) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32584 && (row * 640 + col) <= 32586) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 32587 && (row * 640 + col) <= 32599) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 32600 && (row * 640 + col) <= 32608) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 32609 && (row * 640 + col) <= 32610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32611 && (row * 640 + col) <= 32667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 32668 && (row * 640 + col) <= 32668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32669 && (row * 640 + col) <= 32669) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 32670 && (row * 640 + col) <= 32688) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 32689 && (row * 640 + col) <= 32690) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 32691 && (row * 640 + col) <= 33222) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 33223 && (row * 640 + col) <= 33223) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33224 && (row * 640 + col) <= 33224) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 33225 && (row * 640 + col) <= 33227) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 33228 && (row * 640 + col) <= 33237) color_data <= 12'b111101110010; else
        if ((row * 640 + col) >= 33238 && (row * 640 + col) <= 33247) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 33248 && (row * 640 + col) <= 33249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33250 && (row * 640 + col) <= 33308) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 33309 && (row * 640 + col) <= 33311) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 33312 && (row * 640 + col) <= 33327) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 33328 && (row * 640 + col) <= 33328) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 33329 && (row * 640 + col) <= 33329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33330 && (row * 640 + col) <= 33863) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 33864 && (row * 640 + col) <= 33865) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33866 && (row * 640 + col) <= 33886) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 33887 && (row * 640 + col) <= 33888) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33889 && (row * 640 + col) <= 33950) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 33951 && (row * 640 + col) <= 33952) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33953 && (row * 640 + col) <= 33965) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 33966 && (row * 640 + col) <= 33968) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 33969 && (row * 640 + col) <= 34504) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 34505 && (row * 640 + col) <= 34505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34506 && (row * 640 + col) <= 34506) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 34507 && (row * 640 + col) <= 34525) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 34526 && (row * 640 + col) <= 34527) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34528 && (row * 640 + col) <= 34591) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 34592 && (row * 640 + col) <= 34592) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34593 && (row * 640 + col) <= 34594) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 34595 && (row * 640 + col) <= 34603) color_data <= 12'b101100000000; else
        if ((row * 640 + col) >= 34604 && (row * 640 + col) <= 34604) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 34605 && (row * 640 + col) <= 34606) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 34607 && (row * 640 + col) <= 35145) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 35146 && (row * 640 + col) <= 35148) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35149 && (row * 640 + col) <= 35163) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 35164 && (row * 640 + col) <= 35166) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35167 && (row * 640 + col) <= 35233) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 35234 && (row * 640 + col) <= 35243) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 35244 && (row * 640 + col) <= 35244) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35245 && (row * 640 + col) <= 35787) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 35788 && (row * 640 + col) <= 35789) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35790 && (row * 640 + col) <= 35790) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 35791 && (row * 640 + col) <= 35801) color_data <= 12'b111001110010; else
        if ((row * 640 + col) >= 35802 && (row * 640 + col) <= 35804) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 35805 && (row * 640 + col) <= 35874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 35875 && (row * 640 + col) <= 36429) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 36430 && (row * 640 + col) <= 36430) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36431 && (row * 640 + col) <= 36440) color_data <= 12'b000100000000; else
        if ((row * 640 + col) >= 36441 && (row * 640 + col) <= 36442) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 36443 && (row * 640 + col) <= 36514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 36515 && (row * 640 + col) <= 37082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 37083 && (row * 640 + col) <= 37154) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 37155 && (row * 640 + col) <= 37722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 37723 && (row * 640 + col) <= 37794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 37795 && (row * 640 + col) <= 38362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 38363 && (row * 640 + col) <= 38434) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 38435 && (row * 640 + col) <= 39002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 39003 && (row * 640 + col) <= 39074) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 39075 && (row * 640 + col) <= 39642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 39643 && (row * 640 + col) <= 39714) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 39715 && (row * 640 + col) <= 40282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 40283 && (row * 640 + col) <= 40354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 40355 && (row * 640 + col) <= 40922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 40923 && (row * 640 + col) <= 40994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 40995 && (row * 640 + col) <= 41562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 41563 && (row * 640 + col) <= 41634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 41635 && (row * 640 + col) <= 42202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 42203 && (row * 640 + col) <= 42274) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 42275 && (row * 640 + col) <= 42842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 42843 && (row * 640 + col) <= 42914) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 42915 && (row * 640 + col) <= 43482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 43483 && (row * 640 + col) <= 43554) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 43555 && (row * 640 + col) <= 44122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 44123 && (row * 640 + col) <= 44194) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 44195 && (row * 640 + col) <= 44762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 44763 && (row * 640 + col) <= 44834) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 44835 && (row * 640 + col) <= 45402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 45403 && (row * 640 + col) <= 45474) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 45475 && (row * 640 + col) <= 46042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 46043 && (row * 640 + col) <= 46114) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 46115 && (row * 640 + col) <= 46682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 46683 && (row * 640 + col) <= 46754) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 46755 && (row * 640 + col) <= 47322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 47323 && (row * 640 + col) <= 47394) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 47395 && (row * 640 + col) <= 47962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 47963 && (row * 640 + col) <= 48034) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 48035 && (row * 640 + col) <= 48602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 48603 && (row * 640 + col) <= 48674) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 48675 && (row * 640 + col) <= 49242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 49243 && (row * 640 + col) <= 49314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 49315 && (row * 640 + col) <= 49882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 49883 && (row * 640 + col) <= 49954) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 49955 && (row * 640 + col) <= 50522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 50523 && (row * 640 + col) <= 50594) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 50595 && (row * 640 + col) <= 51162) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 51163 && (row * 640 + col) <= 51234) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 51235 && (row * 640 + col) <= 51802) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 51803 && (row * 640 + col) <= 51874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 51875 && (row * 640 + col) <= 52442) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 52443 && (row * 640 + col) <= 52514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 52515 && (row * 640 + col) <= 53082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 53083 && (row * 640 + col) <= 53154) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 53155 && (row * 640 + col) <= 53722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 53723 && (row * 640 + col) <= 53794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 53795 && (row * 640 + col) <= 54362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 54363 && (row * 640 + col) <= 54434) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 54435 && (row * 640 + col) <= 55002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 55003 && (row * 640 + col) <= 55074) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 55075 && (row * 640 + col) <= 55642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 55643 && (row * 640 + col) <= 55714) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 55715 && (row * 640 + col) <= 56282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56283 && (row * 640 + col) <= 56354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 56355 && (row * 640 + col) <= 56391) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56392 && (row * 640 + col) <= 56426) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56427 && (row * 640 + col) <= 56433) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56434 && (row * 640 + col) <= 56468) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56469 && (row * 640 + col) <= 56475) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56476 && (row * 640 + col) <= 56489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56490 && (row * 640 + col) <= 56496) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56497 && (row * 640 + col) <= 56510) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56511 && (row * 640 + col) <= 56517) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56518 && (row * 640 + col) <= 56545) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56546 && (row * 640 + col) <= 56552) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56553 && (row * 640 + col) <= 56580) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56581 && (row * 640 + col) <= 56601) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56602 && (row * 640 + col) <= 56636) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56637 && (row * 640 + col) <= 56643) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56644 && (row * 640 + col) <= 56678) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56679 && (row * 640 + col) <= 56685) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56686 && (row * 640 + col) <= 56713) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56714 && (row * 640 + col) <= 56720) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56721 && (row * 640 + col) <= 56755) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56756 && (row * 640 + col) <= 56762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56763 && (row * 640 + col) <= 56776) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56777 && (row * 640 + col) <= 56783) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56784 && (row * 640 + col) <= 56797) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56798 && (row * 640 + col) <= 56804) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56805 && (row * 640 + col) <= 56839) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56840 && (row * 640 + col) <= 56846) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56847 && (row * 640 + col) <= 56881) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 56882 && (row * 640 + col) <= 56922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56923 && (row * 640 + col) <= 56994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 56995 && (row * 640 + col) <= 57031) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57032 && (row * 640 + col) <= 57066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57067 && (row * 640 + col) <= 57073) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57074 && (row * 640 + col) <= 57108) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57109 && (row * 640 + col) <= 57115) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57116 && (row * 640 + col) <= 57129) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57130 && (row * 640 + col) <= 57136) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57137 && (row * 640 + col) <= 57150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57151 && (row * 640 + col) <= 57157) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57158 && (row * 640 + col) <= 57185) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57186 && (row * 640 + col) <= 57192) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57193 && (row * 640 + col) <= 57220) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57221 && (row * 640 + col) <= 57241) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57242 && (row * 640 + col) <= 57276) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57277 && (row * 640 + col) <= 57283) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57284 && (row * 640 + col) <= 57318) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57319 && (row * 640 + col) <= 57325) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57326 && (row * 640 + col) <= 57353) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57354 && (row * 640 + col) <= 57360) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57361 && (row * 640 + col) <= 57395) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57396 && (row * 640 + col) <= 57402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57403 && (row * 640 + col) <= 57416) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57417 && (row * 640 + col) <= 57423) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57424 && (row * 640 + col) <= 57437) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57438 && (row * 640 + col) <= 57444) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57445 && (row * 640 + col) <= 57479) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57480 && (row * 640 + col) <= 57486) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57487 && (row * 640 + col) <= 57521) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57522 && (row * 640 + col) <= 57562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57563 && (row * 640 + col) <= 57634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 57635 && (row * 640 + col) <= 57671) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57672 && (row * 640 + col) <= 57706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57707 && (row * 640 + col) <= 57713) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57714 && (row * 640 + col) <= 57748) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57749 && (row * 640 + col) <= 57755) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57756 && (row * 640 + col) <= 57769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57770 && (row * 640 + col) <= 57776) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57777 && (row * 640 + col) <= 57790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57791 && (row * 640 + col) <= 57797) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57798 && (row * 640 + col) <= 57825) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57826 && (row * 640 + col) <= 57832) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57833 && (row * 640 + col) <= 57860) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57861 && (row * 640 + col) <= 57881) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57882 && (row * 640 + col) <= 57916) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57917 && (row * 640 + col) <= 57923) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57924 && (row * 640 + col) <= 57958) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57959 && (row * 640 + col) <= 57965) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57966 && (row * 640 + col) <= 57993) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 57994 && (row * 640 + col) <= 58000) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58001 && (row * 640 + col) <= 58035) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58036 && (row * 640 + col) <= 58042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58043 && (row * 640 + col) <= 58056) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58057 && (row * 640 + col) <= 58063) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58064 && (row * 640 + col) <= 58077) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58078 && (row * 640 + col) <= 58084) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58085 && (row * 640 + col) <= 58119) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58120 && (row * 640 + col) <= 58126) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58127 && (row * 640 + col) <= 58161) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58162 && (row * 640 + col) <= 58202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58203 && (row * 640 + col) <= 58274) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 58275 && (row * 640 + col) <= 58311) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58312 && (row * 640 + col) <= 58346) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58347 && (row * 640 + col) <= 58353) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58354 && (row * 640 + col) <= 58388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58389 && (row * 640 + col) <= 58395) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58396 && (row * 640 + col) <= 58409) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58410 && (row * 640 + col) <= 58416) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58417 && (row * 640 + col) <= 58430) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58431 && (row * 640 + col) <= 58437) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58438 && (row * 640 + col) <= 58465) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58466 && (row * 640 + col) <= 58472) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58473 && (row * 640 + col) <= 58500) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58501 && (row * 640 + col) <= 58521) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58522 && (row * 640 + col) <= 58556) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58557 && (row * 640 + col) <= 58563) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58564 && (row * 640 + col) <= 58598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58599 && (row * 640 + col) <= 58605) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58606 && (row * 640 + col) <= 58633) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58634 && (row * 640 + col) <= 58640) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58641 && (row * 640 + col) <= 58675) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58676 && (row * 640 + col) <= 58682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58683 && (row * 640 + col) <= 58696) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58697 && (row * 640 + col) <= 58703) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58704 && (row * 640 + col) <= 58717) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58718 && (row * 640 + col) <= 58724) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58725 && (row * 640 + col) <= 58759) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58760 && (row * 640 + col) <= 58766) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58767 && (row * 640 + col) <= 58801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58802 && (row * 640 + col) <= 58842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58843 && (row * 640 + col) <= 58914) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 58915 && (row * 640 + col) <= 58951) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58952 && (row * 640 + col) <= 58986) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 58987 && (row * 640 + col) <= 58993) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58994 && (row * 640 + col) <= 59028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59029 && (row * 640 + col) <= 59035) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59036 && (row * 640 + col) <= 59049) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59050 && (row * 640 + col) <= 59056) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59057 && (row * 640 + col) <= 59070) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59071 && (row * 640 + col) <= 59077) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59078 && (row * 640 + col) <= 59105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59106 && (row * 640 + col) <= 59112) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59113 && (row * 640 + col) <= 59140) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59141 && (row * 640 + col) <= 59161) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59162 && (row * 640 + col) <= 59196) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59197 && (row * 640 + col) <= 59203) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59204 && (row * 640 + col) <= 59238) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59239 && (row * 640 + col) <= 59245) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59246 && (row * 640 + col) <= 59273) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59274 && (row * 640 + col) <= 59280) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59281 && (row * 640 + col) <= 59315) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59316 && (row * 640 + col) <= 59322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59323 && (row * 640 + col) <= 59336) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59337 && (row * 640 + col) <= 59343) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59344 && (row * 640 + col) <= 59357) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59358 && (row * 640 + col) <= 59364) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59365 && (row * 640 + col) <= 59399) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59400 && (row * 640 + col) <= 59406) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59407 && (row * 640 + col) <= 59441) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59442 && (row * 640 + col) <= 59482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59483 && (row * 640 + col) <= 59554) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 59555 && (row * 640 + col) <= 59591) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59592 && (row * 640 + col) <= 59626) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59627 && (row * 640 + col) <= 59633) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59634 && (row * 640 + col) <= 59668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59669 && (row * 640 + col) <= 59675) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59676 && (row * 640 + col) <= 59689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59690 && (row * 640 + col) <= 59696) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59697 && (row * 640 + col) <= 59710) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59711 && (row * 640 + col) <= 59717) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59718 && (row * 640 + col) <= 59745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59746 && (row * 640 + col) <= 59752) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59753 && (row * 640 + col) <= 59780) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59781 && (row * 640 + col) <= 59801) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59802 && (row * 640 + col) <= 59836) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59837 && (row * 640 + col) <= 59843) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59844 && (row * 640 + col) <= 59878) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59879 && (row * 640 + col) <= 59885) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59886 && (row * 640 + col) <= 59913) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59914 && (row * 640 + col) <= 59920) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59921 && (row * 640 + col) <= 59955) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59956 && (row * 640 + col) <= 59962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59963 && (row * 640 + col) <= 59976) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59977 && (row * 640 + col) <= 59983) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59984 && (row * 640 + col) <= 59997) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 59998 && (row * 640 + col) <= 60004) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60005 && (row * 640 + col) <= 60039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60040 && (row * 640 + col) <= 60046) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60047 && (row * 640 + col) <= 60081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60082 && (row * 640 + col) <= 60122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60123 && (row * 640 + col) <= 60194) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 60195 && (row * 640 + col) <= 60231) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60232 && (row * 640 + col) <= 60266) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60267 && (row * 640 + col) <= 60273) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60274 && (row * 640 + col) <= 60308) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60309 && (row * 640 + col) <= 60315) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60316 && (row * 640 + col) <= 60329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60330 && (row * 640 + col) <= 60336) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60337 && (row * 640 + col) <= 60350) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60351 && (row * 640 + col) <= 60357) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60358 && (row * 640 + col) <= 60385) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60386 && (row * 640 + col) <= 60392) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60393 && (row * 640 + col) <= 60420) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60421 && (row * 640 + col) <= 60441) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60442 && (row * 640 + col) <= 60476) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60477 && (row * 640 + col) <= 60483) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60484 && (row * 640 + col) <= 60518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60519 && (row * 640 + col) <= 60525) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60526 && (row * 640 + col) <= 60553) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60554 && (row * 640 + col) <= 60560) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60561 && (row * 640 + col) <= 60595) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60596 && (row * 640 + col) <= 60602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60603 && (row * 640 + col) <= 60616) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60617 && (row * 640 + col) <= 60623) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60624 && (row * 640 + col) <= 60637) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60638 && (row * 640 + col) <= 60644) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60645 && (row * 640 + col) <= 60679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60680 && (row * 640 + col) <= 60686) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60687 && (row * 640 + col) <= 60721) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60722 && (row * 640 + col) <= 60762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60763 && (row * 640 + col) <= 60834) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 60835 && (row * 640 + col) <= 60871) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60872 && (row * 640 + col) <= 60885) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60886 && (row * 640 + col) <= 60892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60893 && (row * 640 + col) <= 60906) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60907 && (row * 640 + col) <= 60913) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60914 && (row * 640 + col) <= 60927) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60928 && (row * 640 + col) <= 60934) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60935 && (row * 640 + col) <= 60948) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60949 && (row * 640 + col) <= 60955) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60956 && (row * 640 + col) <= 60969) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60970 && (row * 640 + col) <= 60976) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60977 && (row * 640 + col) <= 60990) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 60991 && (row * 640 + col) <= 61004) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61005 && (row * 640 + col) <= 61018) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61019 && (row * 640 + col) <= 61039) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61040 && (row * 640 + col) <= 61053) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61054 && (row * 640 + col) <= 61081) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61082 && (row * 640 + col) <= 61095) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61096 && (row * 640 + col) <= 61102) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61103 && (row * 640 + col) <= 61116) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61117 && (row * 640 + col) <= 61123) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61124 && (row * 640 + col) <= 61137) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61138 && (row * 640 + col) <= 61144) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61145 && (row * 640 + col) <= 61158) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61159 && (row * 640 + col) <= 61172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61173 && (row * 640 + col) <= 61186) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61187 && (row * 640 + col) <= 61200) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61201 && (row * 640 + col) <= 61214) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61215 && (row * 640 + col) <= 61221) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61222 && (row * 640 + col) <= 61235) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61236 && (row * 640 + col) <= 61242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61243 && (row * 640 + col) <= 61256) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61257 && (row * 640 + col) <= 61263) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61264 && (row * 640 + col) <= 61277) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61278 && (row * 640 + col) <= 61284) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61285 && (row * 640 + col) <= 61298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61299 && (row * 640 + col) <= 61305) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61306 && (row * 640 + col) <= 61319) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61320 && (row * 640 + col) <= 61326) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61327 && (row * 640 + col) <= 61340) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61341 && (row * 640 + col) <= 61347) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61348 && (row * 640 + col) <= 61361) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61362 && (row * 640 + col) <= 61402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61403 && (row * 640 + col) <= 61474) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 61475 && (row * 640 + col) <= 61511) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61512 && (row * 640 + col) <= 61525) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61526 && (row * 640 + col) <= 61532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61533 && (row * 640 + col) <= 61546) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61547 && (row * 640 + col) <= 61553) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61554 && (row * 640 + col) <= 61567) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61568 && (row * 640 + col) <= 61574) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61575 && (row * 640 + col) <= 61588) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61589 && (row * 640 + col) <= 61595) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61596 && (row * 640 + col) <= 61609) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61610 && (row * 640 + col) <= 61616) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61617 && (row * 640 + col) <= 61630) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61631 && (row * 640 + col) <= 61644) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61645 && (row * 640 + col) <= 61658) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61659 && (row * 640 + col) <= 61679) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61680 && (row * 640 + col) <= 61693) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61694 && (row * 640 + col) <= 61721) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61722 && (row * 640 + col) <= 61735) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61736 && (row * 640 + col) <= 61742) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61743 && (row * 640 + col) <= 61756) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61757 && (row * 640 + col) <= 61763) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61764 && (row * 640 + col) <= 61777) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61778 && (row * 640 + col) <= 61784) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61785 && (row * 640 + col) <= 61798) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61799 && (row * 640 + col) <= 61812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61813 && (row * 640 + col) <= 61826) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61827 && (row * 640 + col) <= 61840) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61841 && (row * 640 + col) <= 61854) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61855 && (row * 640 + col) <= 61861) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61862 && (row * 640 + col) <= 61875) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61876 && (row * 640 + col) <= 61882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61883 && (row * 640 + col) <= 61896) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61897 && (row * 640 + col) <= 61903) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61904 && (row * 640 + col) <= 61917) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61918 && (row * 640 + col) <= 61924) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61925 && (row * 640 + col) <= 61938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61939 && (row * 640 + col) <= 61945) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61946 && (row * 640 + col) <= 61959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61960 && (row * 640 + col) <= 61966) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61967 && (row * 640 + col) <= 61980) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 61981 && (row * 640 + col) <= 61987) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61988 && (row * 640 + col) <= 62001) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62002 && (row * 640 + col) <= 62042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62043 && (row * 640 + col) <= 62114) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 62115 && (row * 640 + col) <= 62151) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62152 && (row * 640 + col) <= 62165) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62166 && (row * 640 + col) <= 62172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62173 && (row * 640 + col) <= 62186) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62187 && (row * 640 + col) <= 62193) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62194 && (row * 640 + col) <= 62207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62208 && (row * 640 + col) <= 62214) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62215 && (row * 640 + col) <= 62228) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62229 && (row * 640 + col) <= 62235) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62236 && (row * 640 + col) <= 62249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62250 && (row * 640 + col) <= 62256) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62257 && (row * 640 + col) <= 62270) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62271 && (row * 640 + col) <= 62284) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62285 && (row * 640 + col) <= 62298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62299 && (row * 640 + col) <= 62319) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62320 && (row * 640 + col) <= 62333) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62334 && (row * 640 + col) <= 62361) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62362 && (row * 640 + col) <= 62375) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62376 && (row * 640 + col) <= 62382) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62383 && (row * 640 + col) <= 62396) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62397 && (row * 640 + col) <= 62403) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62404 && (row * 640 + col) <= 62417) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62418 && (row * 640 + col) <= 62424) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62425 && (row * 640 + col) <= 62438) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62439 && (row * 640 + col) <= 62452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62453 && (row * 640 + col) <= 62466) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62467 && (row * 640 + col) <= 62480) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62481 && (row * 640 + col) <= 62494) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62495 && (row * 640 + col) <= 62501) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62502 && (row * 640 + col) <= 62515) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62516 && (row * 640 + col) <= 62522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62523 && (row * 640 + col) <= 62536) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62537 && (row * 640 + col) <= 62543) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62544 && (row * 640 + col) <= 62557) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62558 && (row * 640 + col) <= 62564) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62565 && (row * 640 + col) <= 62578) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62579 && (row * 640 + col) <= 62585) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62586 && (row * 640 + col) <= 62599) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62600 && (row * 640 + col) <= 62606) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62607 && (row * 640 + col) <= 62620) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62621 && (row * 640 + col) <= 62627) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62628 && (row * 640 + col) <= 62641) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62642 && (row * 640 + col) <= 62682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62683 && (row * 640 + col) <= 62754) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 62755 && (row * 640 + col) <= 62791) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62792 && (row * 640 + col) <= 62805) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62806 && (row * 640 + col) <= 62812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62813 && (row * 640 + col) <= 62826) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62827 && (row * 640 + col) <= 62833) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62834 && (row * 640 + col) <= 62847) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62848 && (row * 640 + col) <= 62854) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62855 && (row * 640 + col) <= 62868) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62869 && (row * 640 + col) <= 62875) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62876 && (row * 640 + col) <= 62889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62890 && (row * 640 + col) <= 62896) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62897 && (row * 640 + col) <= 62910) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62911 && (row * 640 + col) <= 62924) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62925 && (row * 640 + col) <= 62938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62939 && (row * 640 + col) <= 62959) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62960 && (row * 640 + col) <= 62973) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 62974 && (row * 640 + col) <= 63001) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63002 && (row * 640 + col) <= 63015) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63016 && (row * 640 + col) <= 63022) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63023 && (row * 640 + col) <= 63036) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63037 && (row * 640 + col) <= 63043) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63044 && (row * 640 + col) <= 63057) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63058 && (row * 640 + col) <= 63064) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63065 && (row * 640 + col) <= 63078) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63079 && (row * 640 + col) <= 63092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63093 && (row * 640 + col) <= 63106) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63107 && (row * 640 + col) <= 63120) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63121 && (row * 640 + col) <= 63134) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63135 && (row * 640 + col) <= 63141) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63142 && (row * 640 + col) <= 63155) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63156 && (row * 640 + col) <= 63162) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63163 && (row * 640 + col) <= 63176) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63177 && (row * 640 + col) <= 63183) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63184 && (row * 640 + col) <= 63197) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63198 && (row * 640 + col) <= 63204) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63205 && (row * 640 + col) <= 63218) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63219 && (row * 640 + col) <= 63225) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63226 && (row * 640 + col) <= 63239) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63240 && (row * 640 + col) <= 63246) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63247 && (row * 640 + col) <= 63260) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63261 && (row * 640 + col) <= 63267) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63268 && (row * 640 + col) <= 63281) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63282 && (row * 640 + col) <= 63322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63323 && (row * 640 + col) <= 63394) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 63395 && (row * 640 + col) <= 63431) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63432 && (row * 640 + col) <= 63445) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63446 && (row * 640 + col) <= 63452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63453 && (row * 640 + col) <= 63466) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63467 && (row * 640 + col) <= 63473) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63474 && (row * 640 + col) <= 63487) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63488 && (row * 640 + col) <= 63494) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63495 && (row * 640 + col) <= 63508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63509 && (row * 640 + col) <= 63515) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63516 && (row * 640 + col) <= 63529) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63530 && (row * 640 + col) <= 63536) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63537 && (row * 640 + col) <= 63550) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63551 && (row * 640 + col) <= 63564) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63565 && (row * 640 + col) <= 63578) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63579 && (row * 640 + col) <= 63599) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63600 && (row * 640 + col) <= 63613) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63614 && (row * 640 + col) <= 63641) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63642 && (row * 640 + col) <= 63655) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63656 && (row * 640 + col) <= 63662) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63663 && (row * 640 + col) <= 63676) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63677 && (row * 640 + col) <= 63683) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63684 && (row * 640 + col) <= 63697) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63698 && (row * 640 + col) <= 63704) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63705 && (row * 640 + col) <= 63718) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63719 && (row * 640 + col) <= 63732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63733 && (row * 640 + col) <= 63746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63747 && (row * 640 + col) <= 63760) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63761 && (row * 640 + col) <= 63774) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63775 && (row * 640 + col) <= 63781) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63782 && (row * 640 + col) <= 63795) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63796 && (row * 640 + col) <= 63802) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63803 && (row * 640 + col) <= 63816) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63817 && (row * 640 + col) <= 63823) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63824 && (row * 640 + col) <= 63837) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63838 && (row * 640 + col) <= 63844) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63845 && (row * 640 + col) <= 63858) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63859 && (row * 640 + col) <= 63865) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63866 && (row * 640 + col) <= 63879) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63880 && (row * 640 + col) <= 63886) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63887 && (row * 640 + col) <= 63900) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63901 && (row * 640 + col) <= 63907) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63908 && (row * 640 + col) <= 63921) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 63922 && (row * 640 + col) <= 63962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63963 && (row * 640 + col) <= 64034) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 64035 && (row * 640 + col) <= 64071) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64072 && (row * 640 + col) <= 64085) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64086 && (row * 640 + col) <= 64092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64093 && (row * 640 + col) <= 64106) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64107 && (row * 640 + col) <= 64113) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64114 && (row * 640 + col) <= 64127) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64128 && (row * 640 + col) <= 64134) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64135 && (row * 640 + col) <= 64148) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64149 && (row * 640 + col) <= 64155) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64156 && (row * 640 + col) <= 64169) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64170 && (row * 640 + col) <= 64176) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64177 && (row * 640 + col) <= 64190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64191 && (row * 640 + col) <= 64204) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64205 && (row * 640 + col) <= 64218) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64219 && (row * 640 + col) <= 64239) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64240 && (row * 640 + col) <= 64253) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64254 && (row * 640 + col) <= 64281) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64282 && (row * 640 + col) <= 64295) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64296 && (row * 640 + col) <= 64302) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64303 && (row * 640 + col) <= 64316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64317 && (row * 640 + col) <= 64323) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64324 && (row * 640 + col) <= 64337) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64338 && (row * 640 + col) <= 64344) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64345 && (row * 640 + col) <= 64358) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64359 && (row * 640 + col) <= 64372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64373 && (row * 640 + col) <= 64386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64387 && (row * 640 + col) <= 64400) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64401 && (row * 640 + col) <= 64414) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64415 && (row * 640 + col) <= 64421) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64422 && (row * 640 + col) <= 64435) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64436 && (row * 640 + col) <= 64442) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64443 && (row * 640 + col) <= 64456) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64457 && (row * 640 + col) <= 64463) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64464 && (row * 640 + col) <= 64477) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64478 && (row * 640 + col) <= 64484) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64485 && (row * 640 + col) <= 64498) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64499 && (row * 640 + col) <= 64505) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64506 && (row * 640 + col) <= 64519) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64520 && (row * 640 + col) <= 64526) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64527 && (row * 640 + col) <= 64540) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64541 && (row * 640 + col) <= 64547) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64548 && (row * 640 + col) <= 64561) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64562 && (row * 640 + col) <= 64602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64603 && (row * 640 + col) <= 64674) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 64675 && (row * 640 + col) <= 64711) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64712 && (row * 640 + col) <= 64725) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64726 && (row * 640 + col) <= 64732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64733 && (row * 640 + col) <= 64746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64747 && (row * 640 + col) <= 64753) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64754 && (row * 640 + col) <= 64767) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64768 && (row * 640 + col) <= 64774) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64775 && (row * 640 + col) <= 64788) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64789 && (row * 640 + col) <= 64795) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64796 && (row * 640 + col) <= 64809) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64810 && (row * 640 + col) <= 64816) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64817 && (row * 640 + col) <= 64830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64831 && (row * 640 + col) <= 64844) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64845 && (row * 640 + col) <= 64858) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64859 && (row * 640 + col) <= 64879) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64880 && (row * 640 + col) <= 64893) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64894 && (row * 640 + col) <= 64921) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64922 && (row * 640 + col) <= 64935) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64936 && (row * 640 + col) <= 64942) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64943 && (row * 640 + col) <= 64956) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64957 && (row * 640 + col) <= 64963) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64964 && (row * 640 + col) <= 64977) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64978 && (row * 640 + col) <= 64984) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64985 && (row * 640 + col) <= 64998) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 64999 && (row * 640 + col) <= 65012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65013 && (row * 640 + col) <= 65026) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65027 && (row * 640 + col) <= 65040) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65041 && (row * 640 + col) <= 65054) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65055 && (row * 640 + col) <= 65061) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65062 && (row * 640 + col) <= 65075) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65076 && (row * 640 + col) <= 65082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65083 && (row * 640 + col) <= 65096) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65097 && (row * 640 + col) <= 65103) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65104 && (row * 640 + col) <= 65117) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65118 && (row * 640 + col) <= 65124) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65125 && (row * 640 + col) <= 65138) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65139 && (row * 640 + col) <= 65145) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65146 && (row * 640 + col) <= 65159) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65160 && (row * 640 + col) <= 65166) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65167 && (row * 640 + col) <= 65180) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65181 && (row * 640 + col) <= 65187) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65188 && (row * 640 + col) <= 65201) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65202 && (row * 640 + col) <= 65242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65243 && (row * 640 + col) <= 65314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 65315 && (row * 640 + col) <= 65351) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65352 && (row * 640 + col) <= 65365) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65366 && (row * 640 + col) <= 65393) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65394 && (row * 640 + col) <= 65407) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65408 && (row * 640 + col) <= 65414) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65415 && (row * 640 + col) <= 65428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65429 && (row * 640 + col) <= 65435) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65436 && (row * 640 + col) <= 65449) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65450 && (row * 640 + col) <= 65456) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65457 && (row * 640 + col) <= 65470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65471 && (row * 640 + col) <= 65484) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65485 && (row * 640 + col) <= 65498) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65499 && (row * 640 + col) <= 65519) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65520 && (row * 640 + col) <= 65533) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65534 && (row * 640 + col) <= 65561) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65562 && (row * 640 + col) <= 65575) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65576 && (row * 640 + col) <= 65603) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65604 && (row * 640 + col) <= 65617) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65618 && (row * 640 + col) <= 65624) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65625 && (row * 640 + col) <= 65638) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65639 && (row * 640 + col) <= 65652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65653 && (row * 640 + col) <= 65666) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65667 && (row * 640 + col) <= 65680) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65681 && (row * 640 + col) <= 65694) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65695 && (row * 640 + col) <= 65722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65723 && (row * 640 + col) <= 65736) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65737 && (row * 640 + col) <= 65743) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65744 && (row * 640 + col) <= 65757) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65758 && (row * 640 + col) <= 65764) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65765 && (row * 640 + col) <= 65778) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65779 && (row * 640 + col) <= 65806) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65807 && (row * 640 + col) <= 65820) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65821 && (row * 640 + col) <= 65827) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65828 && (row * 640 + col) <= 65841) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 65842 && (row * 640 + col) <= 65882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65883 && (row * 640 + col) <= 65954) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 65955 && (row * 640 + col) <= 65991) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65992 && (row * 640 + col) <= 66005) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66006 && (row * 640 + col) <= 66033) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66034 && (row * 640 + col) <= 66047) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66048 && (row * 640 + col) <= 66054) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66055 && (row * 640 + col) <= 66068) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66069 && (row * 640 + col) <= 66075) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66076 && (row * 640 + col) <= 66089) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66090 && (row * 640 + col) <= 66096) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66097 && (row * 640 + col) <= 66110) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66111 && (row * 640 + col) <= 66124) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66125 && (row * 640 + col) <= 66138) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66139 && (row * 640 + col) <= 66159) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66160 && (row * 640 + col) <= 66173) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66174 && (row * 640 + col) <= 66201) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66202 && (row * 640 + col) <= 66215) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66216 && (row * 640 + col) <= 66243) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66244 && (row * 640 + col) <= 66257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66258 && (row * 640 + col) <= 66264) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66265 && (row * 640 + col) <= 66278) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66279 && (row * 640 + col) <= 66292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66293 && (row * 640 + col) <= 66306) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66307 && (row * 640 + col) <= 66320) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66321 && (row * 640 + col) <= 66334) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66335 && (row * 640 + col) <= 66362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66363 && (row * 640 + col) <= 66376) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66377 && (row * 640 + col) <= 66383) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66384 && (row * 640 + col) <= 66397) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66398 && (row * 640 + col) <= 66404) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66405 && (row * 640 + col) <= 66418) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66419 && (row * 640 + col) <= 66446) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66447 && (row * 640 + col) <= 66460) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66461 && (row * 640 + col) <= 66467) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66468 && (row * 640 + col) <= 66481) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66482 && (row * 640 + col) <= 66522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66523 && (row * 640 + col) <= 66594) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 66595 && (row * 640 + col) <= 66631) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66632 && (row * 640 + col) <= 66645) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66646 && (row * 640 + col) <= 66673) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66674 && (row * 640 + col) <= 66687) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66688 && (row * 640 + col) <= 66694) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66695 && (row * 640 + col) <= 66708) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66709 && (row * 640 + col) <= 66715) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66716 && (row * 640 + col) <= 66729) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66730 && (row * 640 + col) <= 66736) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66737 && (row * 640 + col) <= 66750) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66751 && (row * 640 + col) <= 66764) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66765 && (row * 640 + col) <= 66778) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66779 && (row * 640 + col) <= 66799) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66800 && (row * 640 + col) <= 66813) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66814 && (row * 640 + col) <= 66841) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66842 && (row * 640 + col) <= 66855) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66856 && (row * 640 + col) <= 66883) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66884 && (row * 640 + col) <= 66897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66898 && (row * 640 + col) <= 66904) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66905 && (row * 640 + col) <= 66918) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66919 && (row * 640 + col) <= 66932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66933 && (row * 640 + col) <= 66946) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66947 && (row * 640 + col) <= 66960) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66961 && (row * 640 + col) <= 66974) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 66975 && (row * 640 + col) <= 67002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67003 && (row * 640 + col) <= 67016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67017 && (row * 640 + col) <= 67023) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67024 && (row * 640 + col) <= 67037) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67038 && (row * 640 + col) <= 67044) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67045 && (row * 640 + col) <= 67058) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67059 && (row * 640 + col) <= 67086) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67087 && (row * 640 + col) <= 67100) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67101 && (row * 640 + col) <= 67107) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67108 && (row * 640 + col) <= 67121) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67122 && (row * 640 + col) <= 67162) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67163 && (row * 640 + col) <= 67234) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 67235 && (row * 640 + col) <= 67271) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67272 && (row * 640 + col) <= 67285) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67286 && (row * 640 + col) <= 67313) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67314 && (row * 640 + col) <= 67327) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67328 && (row * 640 + col) <= 67334) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67335 && (row * 640 + col) <= 67348) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67349 && (row * 640 + col) <= 67355) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67356 && (row * 640 + col) <= 67369) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67370 && (row * 640 + col) <= 67376) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67377 && (row * 640 + col) <= 67390) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67391 && (row * 640 + col) <= 67404) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67405 && (row * 640 + col) <= 67418) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67419 && (row * 640 + col) <= 67439) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67440 && (row * 640 + col) <= 67453) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67454 && (row * 640 + col) <= 67481) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67482 && (row * 640 + col) <= 67495) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67496 && (row * 640 + col) <= 67523) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67524 && (row * 640 + col) <= 67537) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67538 && (row * 640 + col) <= 67544) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67545 && (row * 640 + col) <= 67558) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67559 && (row * 640 + col) <= 67572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67573 && (row * 640 + col) <= 67586) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67587 && (row * 640 + col) <= 67600) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67601 && (row * 640 + col) <= 67614) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67615 && (row * 640 + col) <= 67642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67643 && (row * 640 + col) <= 67656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67657 && (row * 640 + col) <= 67663) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67664 && (row * 640 + col) <= 67677) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67678 && (row * 640 + col) <= 67684) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67685 && (row * 640 + col) <= 67698) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67699 && (row * 640 + col) <= 67726) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67727 && (row * 640 + col) <= 67740) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67741 && (row * 640 + col) <= 67747) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67748 && (row * 640 + col) <= 67761) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67762 && (row * 640 + col) <= 67802) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67803 && (row * 640 + col) <= 67874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 67875 && (row * 640 + col) <= 67911) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67912 && (row * 640 + col) <= 67925) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67926 && (row * 640 + col) <= 67953) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67954 && (row * 640 + col) <= 67967) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67968 && (row * 640 + col) <= 67974) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67975 && (row * 640 + col) <= 67988) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 67989 && (row * 640 + col) <= 67995) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67996 && (row * 640 + col) <= 68009) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68010 && (row * 640 + col) <= 68016) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68017 && (row * 640 + col) <= 68030) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68031 && (row * 640 + col) <= 68044) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68045 && (row * 640 + col) <= 68058) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68059 && (row * 640 + col) <= 68079) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68080 && (row * 640 + col) <= 68093) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68094 && (row * 640 + col) <= 68121) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68122 && (row * 640 + col) <= 68135) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68136 && (row * 640 + col) <= 68163) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68164 && (row * 640 + col) <= 68177) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68178 && (row * 640 + col) <= 68184) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68185 && (row * 640 + col) <= 68198) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68199 && (row * 640 + col) <= 68212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68213 && (row * 640 + col) <= 68226) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68227 && (row * 640 + col) <= 68240) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68241 && (row * 640 + col) <= 68254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68255 && (row * 640 + col) <= 68282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68283 && (row * 640 + col) <= 68296) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68297 && (row * 640 + col) <= 68303) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68304 && (row * 640 + col) <= 68317) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68318 && (row * 640 + col) <= 68324) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68325 && (row * 640 + col) <= 68338) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68339 && (row * 640 + col) <= 68366) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68367 && (row * 640 + col) <= 68380) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68381 && (row * 640 + col) <= 68387) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68388 && (row * 640 + col) <= 68401) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68402 && (row * 640 + col) <= 68442) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68443 && (row * 640 + col) <= 68514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 68515 && (row * 640 + col) <= 68551) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68552 && (row * 640 + col) <= 68565) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68566 && (row * 640 + col) <= 68593) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68594 && (row * 640 + col) <= 68607) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68608 && (row * 640 + col) <= 68614) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68615 && (row * 640 + col) <= 68628) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68629 && (row * 640 + col) <= 68635) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68636 && (row * 640 + col) <= 68649) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68650 && (row * 640 + col) <= 68656) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68657 && (row * 640 + col) <= 68670) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68671 && (row * 640 + col) <= 68684) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68685 && (row * 640 + col) <= 68698) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68699 && (row * 640 + col) <= 68719) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68720 && (row * 640 + col) <= 68733) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68734 && (row * 640 + col) <= 68761) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68762 && (row * 640 + col) <= 68775) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68776 && (row * 640 + col) <= 68803) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68804 && (row * 640 + col) <= 68817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68818 && (row * 640 + col) <= 68824) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68825 && (row * 640 + col) <= 68838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68839 && (row * 640 + col) <= 68852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68853 && (row * 640 + col) <= 68866) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68867 && (row * 640 + col) <= 68880) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68881 && (row * 640 + col) <= 68894) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68895 && (row * 640 + col) <= 68922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68923 && (row * 640 + col) <= 68936) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68937 && (row * 640 + col) <= 68943) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68944 && (row * 640 + col) <= 68957) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68958 && (row * 640 + col) <= 68964) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68965 && (row * 640 + col) <= 68978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 68979 && (row * 640 + col) <= 69006) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69007 && (row * 640 + col) <= 69020) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69021 && (row * 640 + col) <= 69027) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69028 && (row * 640 + col) <= 69041) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69042 && (row * 640 + col) <= 69082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69083 && (row * 640 + col) <= 69154) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 69155 && (row * 640 + col) <= 69191) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69192 && (row * 640 + col) <= 69205) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69206 && (row * 640 + col) <= 69233) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69234 && (row * 640 + col) <= 69247) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69248 && (row * 640 + col) <= 69254) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69255 && (row * 640 + col) <= 69268) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69269 && (row * 640 + col) <= 69275) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69276 && (row * 640 + col) <= 69289) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69290 && (row * 640 + col) <= 69296) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69297 && (row * 640 + col) <= 69310) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69311 && (row * 640 + col) <= 69324) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69325 && (row * 640 + col) <= 69338) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69339 && (row * 640 + col) <= 69359) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69360 && (row * 640 + col) <= 69373) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69374 && (row * 640 + col) <= 69401) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69402 && (row * 640 + col) <= 69415) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69416 && (row * 640 + col) <= 69443) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69444 && (row * 640 + col) <= 69457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69458 && (row * 640 + col) <= 69464) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69465 && (row * 640 + col) <= 69478) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69479 && (row * 640 + col) <= 69492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69493 && (row * 640 + col) <= 69506) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69507 && (row * 640 + col) <= 69520) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69521 && (row * 640 + col) <= 69534) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69535 && (row * 640 + col) <= 69562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69563 && (row * 640 + col) <= 69576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69577 && (row * 640 + col) <= 69583) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69584 && (row * 640 + col) <= 69597) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69598 && (row * 640 + col) <= 69604) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69605 && (row * 640 + col) <= 69618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69619 && (row * 640 + col) <= 69646) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69647 && (row * 640 + col) <= 69660) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69661 && (row * 640 + col) <= 69667) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69668 && (row * 640 + col) <= 69681) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69682 && (row * 640 + col) <= 69722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69723 && (row * 640 + col) <= 69794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 69795 && (row * 640 + col) <= 69831) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69832 && (row * 640 + col) <= 69859) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69860 && (row * 640 + col) <= 69873) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69874 && (row * 640 + col) <= 69901) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69902 && (row * 640 + col) <= 69915) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69916 && (row * 640 + col) <= 69929) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69930 && (row * 640 + col) <= 69936) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69937 && (row * 640 + col) <= 69950) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69951 && (row * 640 + col) <= 69964) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69965 && (row * 640 + col) <= 69978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 69979 && (row * 640 + col) <= 69999) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70000 && (row * 640 + col) <= 70013) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70014 && (row * 640 + col) <= 70041) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70042 && (row * 640 + col) <= 70055) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70056 && (row * 640 + col) <= 70083) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70084 && (row * 640 + col) <= 70118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70119 && (row * 640 + col) <= 70132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70133 && (row * 640 + col) <= 70146) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70147 && (row * 640 + col) <= 70160) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70161 && (row * 640 + col) <= 70174) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70175 && (row * 640 + col) <= 70202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70203 && (row * 640 + col) <= 70237) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70238 && (row * 640 + col) <= 70244) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70245 && (row * 640 + col) <= 70272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70273 && (row * 640 + col) <= 70286) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70287 && (row * 640 + col) <= 70314) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70315 && (row * 640 + col) <= 70362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70363 && (row * 640 + col) <= 70434) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 70435 && (row * 640 + col) <= 70471) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70472 && (row * 640 + col) <= 70499) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70500 && (row * 640 + col) <= 70513) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70514 && (row * 640 + col) <= 70541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70542 && (row * 640 + col) <= 70555) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70556 && (row * 640 + col) <= 70569) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70570 && (row * 640 + col) <= 70576) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70577 && (row * 640 + col) <= 70590) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70591 && (row * 640 + col) <= 70604) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70605 && (row * 640 + col) <= 70618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70619 && (row * 640 + col) <= 70639) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70640 && (row * 640 + col) <= 70653) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70654 && (row * 640 + col) <= 70681) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70682 && (row * 640 + col) <= 70695) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70696 && (row * 640 + col) <= 70723) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70724 && (row * 640 + col) <= 70758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70759 && (row * 640 + col) <= 70772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70773 && (row * 640 + col) <= 70786) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70787 && (row * 640 + col) <= 70800) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70801 && (row * 640 + col) <= 70814) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70815 && (row * 640 + col) <= 70842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70843 && (row * 640 + col) <= 70877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70878 && (row * 640 + col) <= 70884) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70885 && (row * 640 + col) <= 70912) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70913 && (row * 640 + col) <= 70926) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70927 && (row * 640 + col) <= 70954) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 70955 && (row * 640 + col) <= 71002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71003 && (row * 640 + col) <= 71074) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 71075 && (row * 640 + col) <= 71111) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71112 && (row * 640 + col) <= 71139) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71140 && (row * 640 + col) <= 71153) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71154 && (row * 640 + col) <= 71181) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71182 && (row * 640 + col) <= 71195) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71196 && (row * 640 + col) <= 71209) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71210 && (row * 640 + col) <= 71216) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71217 && (row * 640 + col) <= 71230) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71231 && (row * 640 + col) <= 71244) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71245 && (row * 640 + col) <= 71258) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71259 && (row * 640 + col) <= 71279) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71280 && (row * 640 + col) <= 71293) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71294 && (row * 640 + col) <= 71321) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71322 && (row * 640 + col) <= 71335) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71336 && (row * 640 + col) <= 71363) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71364 && (row * 640 + col) <= 71398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71399 && (row * 640 + col) <= 71412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71413 && (row * 640 + col) <= 71426) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71427 && (row * 640 + col) <= 71440) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71441 && (row * 640 + col) <= 71454) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71455 && (row * 640 + col) <= 71482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71483 && (row * 640 + col) <= 71517) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71518 && (row * 640 + col) <= 71524) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71525 && (row * 640 + col) <= 71552) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71553 && (row * 640 + col) <= 71566) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71567 && (row * 640 + col) <= 71594) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71595 && (row * 640 + col) <= 71642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71643 && (row * 640 + col) <= 71714) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 71715 && (row * 640 + col) <= 71751) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71752 && (row * 640 + col) <= 71779) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71780 && (row * 640 + col) <= 71793) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71794 && (row * 640 + col) <= 71821) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71822 && (row * 640 + col) <= 71835) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71836 && (row * 640 + col) <= 71849) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71850 && (row * 640 + col) <= 71856) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71857 && (row * 640 + col) <= 71870) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71871 && (row * 640 + col) <= 71884) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71885 && (row * 640 + col) <= 71898) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71899 && (row * 640 + col) <= 71919) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71920 && (row * 640 + col) <= 71933) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71934 && (row * 640 + col) <= 71961) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71962 && (row * 640 + col) <= 71975) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 71976 && (row * 640 + col) <= 72003) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72004 && (row * 640 + col) <= 72038) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72039 && (row * 640 + col) <= 72052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72053 && (row * 640 + col) <= 72066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72067 && (row * 640 + col) <= 72080) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72081 && (row * 640 + col) <= 72094) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72095 && (row * 640 + col) <= 72122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72123 && (row * 640 + col) <= 72157) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72158 && (row * 640 + col) <= 72164) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72165 && (row * 640 + col) <= 72192) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72193 && (row * 640 + col) <= 72206) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72207 && (row * 640 + col) <= 72234) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72235 && (row * 640 + col) <= 72282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72283 && (row * 640 + col) <= 72354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 72355 && (row * 640 + col) <= 72391) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72392 && (row * 640 + col) <= 72419) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72420 && (row * 640 + col) <= 72433) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72434 && (row * 640 + col) <= 72461) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72462 && (row * 640 + col) <= 72475) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72476 && (row * 640 + col) <= 72489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72490 && (row * 640 + col) <= 72496) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72497 && (row * 640 + col) <= 72510) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72511 && (row * 640 + col) <= 72524) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72525 && (row * 640 + col) <= 72538) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72539 && (row * 640 + col) <= 72559) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72560 && (row * 640 + col) <= 72573) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72574 && (row * 640 + col) <= 72601) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72602 && (row * 640 + col) <= 72615) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72616 && (row * 640 + col) <= 72643) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72644 && (row * 640 + col) <= 72678) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72679 && (row * 640 + col) <= 72692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72693 && (row * 640 + col) <= 72706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72707 && (row * 640 + col) <= 72720) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72721 && (row * 640 + col) <= 72734) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72735 && (row * 640 + col) <= 72762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72763 && (row * 640 + col) <= 72797) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72798 && (row * 640 + col) <= 72804) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72805 && (row * 640 + col) <= 72832) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72833 && (row * 640 + col) <= 72846) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72847 && (row * 640 + col) <= 72874) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 72875 && (row * 640 + col) <= 72922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72923 && (row * 640 + col) <= 72994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 72995 && (row * 640 + col) <= 73031) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73032 && (row * 640 + col) <= 73059) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73060 && (row * 640 + col) <= 73073) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73074 && (row * 640 + col) <= 73101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73102 && (row * 640 + col) <= 73115) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73116 && (row * 640 + col) <= 73129) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73130 && (row * 640 + col) <= 73136) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73137 && (row * 640 + col) <= 73150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73151 && (row * 640 + col) <= 73164) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73165 && (row * 640 + col) <= 73178) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73179 && (row * 640 + col) <= 73199) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73200 && (row * 640 + col) <= 73213) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73214 && (row * 640 + col) <= 73241) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73242 && (row * 640 + col) <= 73255) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73256 && (row * 640 + col) <= 73283) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73284 && (row * 640 + col) <= 73318) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73319 && (row * 640 + col) <= 73332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73333 && (row * 640 + col) <= 73346) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73347 && (row * 640 + col) <= 73360) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73361 && (row * 640 + col) <= 73374) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73375 && (row * 640 + col) <= 73402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73403 && (row * 640 + col) <= 73437) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73438 && (row * 640 + col) <= 73444) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73445 && (row * 640 + col) <= 73472) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73473 && (row * 640 + col) <= 73486) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73487 && (row * 640 + col) <= 73514) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73515 && (row * 640 + col) <= 73562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73563 && (row * 640 + col) <= 73634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 73635 && (row * 640 + col) <= 73671) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73672 && (row * 640 + col) <= 73699) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73700 && (row * 640 + col) <= 73713) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73714 && (row * 640 + col) <= 73741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73742 && (row * 640 + col) <= 73755) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73756 && (row * 640 + col) <= 73769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73770 && (row * 640 + col) <= 73776) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73777 && (row * 640 + col) <= 73790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73791 && (row * 640 + col) <= 73804) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73805 && (row * 640 + col) <= 73818) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73819 && (row * 640 + col) <= 73839) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73840 && (row * 640 + col) <= 73853) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73854 && (row * 640 + col) <= 73881) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73882 && (row * 640 + col) <= 73895) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73896 && (row * 640 + col) <= 73923) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73924 && (row * 640 + col) <= 73958) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73959 && (row * 640 + col) <= 73972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73973 && (row * 640 + col) <= 73986) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 73987 && (row * 640 + col) <= 74000) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74001 && (row * 640 + col) <= 74014) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74015 && (row * 640 + col) <= 74042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74043 && (row * 640 + col) <= 74077) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74078 && (row * 640 + col) <= 74084) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74085 && (row * 640 + col) <= 74112) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74113 && (row * 640 + col) <= 74126) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74127 && (row * 640 + col) <= 74154) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74155 && (row * 640 + col) <= 74202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74203 && (row * 640 + col) <= 74274) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 74275 && (row * 640 + col) <= 74311) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74312 && (row * 640 + col) <= 74325) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74326 && (row * 640 + col) <= 74353) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74354 && (row * 640 + col) <= 74367) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74368 && (row * 640 + col) <= 74374) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74375 && (row * 640 + col) <= 74388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74389 && (row * 640 + col) <= 74395) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74396 && (row * 640 + col) <= 74409) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74410 && (row * 640 + col) <= 74416) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74417 && (row * 640 + col) <= 74430) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74431 && (row * 640 + col) <= 74444) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74445 && (row * 640 + col) <= 74458) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74459 && (row * 640 + col) <= 74479) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74480 && (row * 640 + col) <= 74493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74494 && (row * 640 + col) <= 74521) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74522 && (row * 640 + col) <= 74535) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74536 && (row * 640 + col) <= 74563) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74564 && (row * 640 + col) <= 74577) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74578 && (row * 640 + col) <= 74584) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74585 && (row * 640 + col) <= 74598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74599 && (row * 640 + col) <= 74612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74613 && (row * 640 + col) <= 74626) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74627 && (row * 640 + col) <= 74640) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74641 && (row * 640 + col) <= 74654) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74655 && (row * 640 + col) <= 74682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74683 && (row * 640 + col) <= 74696) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74697 && (row * 640 + col) <= 74703) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74704 && (row * 640 + col) <= 74717) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74718 && (row * 640 + col) <= 74724) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74725 && (row * 640 + col) <= 74738) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74739 && (row * 640 + col) <= 74766) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74767 && (row * 640 + col) <= 74780) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74781 && (row * 640 + col) <= 74787) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74788 && (row * 640 + col) <= 74801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74802 && (row * 640 + col) <= 74842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74843 && (row * 640 + col) <= 74914) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 74915 && (row * 640 + col) <= 74951) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74952 && (row * 640 + col) <= 74965) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 74966 && (row * 640 + col) <= 74993) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74994 && (row * 640 + col) <= 75007) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75008 && (row * 640 + col) <= 75014) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75015 && (row * 640 + col) <= 75028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75029 && (row * 640 + col) <= 75035) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75036 && (row * 640 + col) <= 75049) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75050 && (row * 640 + col) <= 75056) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75057 && (row * 640 + col) <= 75070) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75071 && (row * 640 + col) <= 75084) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75085 && (row * 640 + col) <= 75098) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75099 && (row * 640 + col) <= 75119) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75120 && (row * 640 + col) <= 75133) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75134 && (row * 640 + col) <= 75161) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75162 && (row * 640 + col) <= 75175) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75176 && (row * 640 + col) <= 75203) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75204 && (row * 640 + col) <= 75217) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75218 && (row * 640 + col) <= 75224) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75225 && (row * 640 + col) <= 75238) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75239 && (row * 640 + col) <= 75252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75253 && (row * 640 + col) <= 75266) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75267 && (row * 640 + col) <= 75280) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75281 && (row * 640 + col) <= 75294) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75295 && (row * 640 + col) <= 75322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75323 && (row * 640 + col) <= 75336) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75337 && (row * 640 + col) <= 75343) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75344 && (row * 640 + col) <= 75357) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75358 && (row * 640 + col) <= 75364) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75365 && (row * 640 + col) <= 75378) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75379 && (row * 640 + col) <= 75406) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75407 && (row * 640 + col) <= 75420) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75421 && (row * 640 + col) <= 75427) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75428 && (row * 640 + col) <= 75441) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75442 && (row * 640 + col) <= 75482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75483 && (row * 640 + col) <= 75554) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 75555 && (row * 640 + col) <= 75591) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75592 && (row * 640 + col) <= 75605) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75606 && (row * 640 + col) <= 75633) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75634 && (row * 640 + col) <= 75647) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75648 && (row * 640 + col) <= 75654) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75655 && (row * 640 + col) <= 75668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75669 && (row * 640 + col) <= 75675) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75676 && (row * 640 + col) <= 75689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75690 && (row * 640 + col) <= 75696) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75697 && (row * 640 + col) <= 75710) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75711 && (row * 640 + col) <= 75724) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75725 && (row * 640 + col) <= 75738) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75739 && (row * 640 + col) <= 75759) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75760 && (row * 640 + col) <= 75773) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75774 && (row * 640 + col) <= 75801) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75802 && (row * 640 + col) <= 75815) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75816 && (row * 640 + col) <= 75843) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75844 && (row * 640 + col) <= 75857) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75858 && (row * 640 + col) <= 75864) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75865 && (row * 640 + col) <= 75878) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75879 && (row * 640 + col) <= 75892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75893 && (row * 640 + col) <= 75906) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75907 && (row * 640 + col) <= 75920) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75921 && (row * 640 + col) <= 75934) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75935 && (row * 640 + col) <= 75962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75963 && (row * 640 + col) <= 75976) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75977 && (row * 640 + col) <= 75983) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75984 && (row * 640 + col) <= 75997) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 75998 && (row * 640 + col) <= 76004) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76005 && (row * 640 + col) <= 76018) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76019 && (row * 640 + col) <= 76046) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76047 && (row * 640 + col) <= 76060) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76061 && (row * 640 + col) <= 76067) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76068 && (row * 640 + col) <= 76081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76082 && (row * 640 + col) <= 76122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76123 && (row * 640 + col) <= 76194) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 76195 && (row * 640 + col) <= 76231) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76232 && (row * 640 + col) <= 76245) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76246 && (row * 640 + col) <= 76273) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76274 && (row * 640 + col) <= 76287) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76288 && (row * 640 + col) <= 76294) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76295 && (row * 640 + col) <= 76308) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76309 && (row * 640 + col) <= 76315) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76316 && (row * 640 + col) <= 76329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76330 && (row * 640 + col) <= 76336) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76337 && (row * 640 + col) <= 76350) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76351 && (row * 640 + col) <= 76364) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76365 && (row * 640 + col) <= 76378) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76379 && (row * 640 + col) <= 76399) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76400 && (row * 640 + col) <= 76413) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76414 && (row * 640 + col) <= 76441) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76442 && (row * 640 + col) <= 76455) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76456 && (row * 640 + col) <= 76483) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76484 && (row * 640 + col) <= 76497) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76498 && (row * 640 + col) <= 76504) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76505 && (row * 640 + col) <= 76518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76519 && (row * 640 + col) <= 76532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76533 && (row * 640 + col) <= 76546) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76547 && (row * 640 + col) <= 76560) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76561 && (row * 640 + col) <= 76574) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76575 && (row * 640 + col) <= 76602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76603 && (row * 640 + col) <= 76616) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76617 && (row * 640 + col) <= 76623) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76624 && (row * 640 + col) <= 76637) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76638 && (row * 640 + col) <= 76644) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76645 && (row * 640 + col) <= 76658) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76659 && (row * 640 + col) <= 76686) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76687 && (row * 640 + col) <= 76700) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76701 && (row * 640 + col) <= 76707) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76708 && (row * 640 + col) <= 76721) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76722 && (row * 640 + col) <= 76762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76763 && (row * 640 + col) <= 76834) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 76835 && (row * 640 + col) <= 76871) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76872 && (row * 640 + col) <= 76885) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76886 && (row * 640 + col) <= 76913) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76914 && (row * 640 + col) <= 76927) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76928 && (row * 640 + col) <= 76934) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76935 && (row * 640 + col) <= 76948) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76949 && (row * 640 + col) <= 76955) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76956 && (row * 640 + col) <= 76969) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76970 && (row * 640 + col) <= 76976) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76977 && (row * 640 + col) <= 76990) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 76991 && (row * 640 + col) <= 77004) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77005 && (row * 640 + col) <= 77018) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77019 && (row * 640 + col) <= 77039) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77040 && (row * 640 + col) <= 77053) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77054 && (row * 640 + col) <= 77081) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77082 && (row * 640 + col) <= 77095) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77096 && (row * 640 + col) <= 77123) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77124 && (row * 640 + col) <= 77137) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77138 && (row * 640 + col) <= 77144) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77145 && (row * 640 + col) <= 77158) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77159 && (row * 640 + col) <= 77172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77173 && (row * 640 + col) <= 77186) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77187 && (row * 640 + col) <= 77200) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77201 && (row * 640 + col) <= 77214) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77215 && (row * 640 + col) <= 77242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77243 && (row * 640 + col) <= 77256) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77257 && (row * 640 + col) <= 77263) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77264 && (row * 640 + col) <= 77277) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77278 && (row * 640 + col) <= 77284) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77285 && (row * 640 + col) <= 77298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77299 && (row * 640 + col) <= 77326) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77327 && (row * 640 + col) <= 77340) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77341 && (row * 640 + col) <= 77347) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77348 && (row * 640 + col) <= 77361) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77362 && (row * 640 + col) <= 77402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77403 && (row * 640 + col) <= 77474) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 77475 && (row * 640 + col) <= 77511) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77512 && (row * 640 + col) <= 77525) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77526 && (row * 640 + col) <= 77553) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77554 && (row * 640 + col) <= 77567) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77568 && (row * 640 + col) <= 77574) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77575 && (row * 640 + col) <= 77588) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77589 && (row * 640 + col) <= 77595) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77596 && (row * 640 + col) <= 77609) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77610 && (row * 640 + col) <= 77616) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77617 && (row * 640 + col) <= 77630) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77631 && (row * 640 + col) <= 77644) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77645 && (row * 640 + col) <= 77658) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77659 && (row * 640 + col) <= 77679) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77680 && (row * 640 + col) <= 77693) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77694 && (row * 640 + col) <= 77721) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77722 && (row * 640 + col) <= 77735) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77736 && (row * 640 + col) <= 77763) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77764 && (row * 640 + col) <= 77777) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77778 && (row * 640 + col) <= 77784) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77785 && (row * 640 + col) <= 77798) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77799 && (row * 640 + col) <= 77812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77813 && (row * 640 + col) <= 77826) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77827 && (row * 640 + col) <= 77840) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77841 && (row * 640 + col) <= 77854) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77855 && (row * 640 + col) <= 77882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77883 && (row * 640 + col) <= 77896) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77897 && (row * 640 + col) <= 77903) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77904 && (row * 640 + col) <= 77917) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77918 && (row * 640 + col) <= 77924) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77925 && (row * 640 + col) <= 77938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77939 && (row * 640 + col) <= 77966) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77967 && (row * 640 + col) <= 77980) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 77981 && (row * 640 + col) <= 77987) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77988 && (row * 640 + col) <= 78001) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78002 && (row * 640 + col) <= 78042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78043 && (row * 640 + col) <= 78114) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 78115 && (row * 640 + col) <= 78151) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78152 && (row * 640 + col) <= 78165) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78166 && (row * 640 + col) <= 78193) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78194 && (row * 640 + col) <= 78207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78208 && (row * 640 + col) <= 78214) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78215 && (row * 640 + col) <= 78228) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78229 && (row * 640 + col) <= 78235) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78236 && (row * 640 + col) <= 78249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78250 && (row * 640 + col) <= 78256) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78257 && (row * 640 + col) <= 78270) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78271 && (row * 640 + col) <= 78284) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78285 && (row * 640 + col) <= 78298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78299 && (row * 640 + col) <= 78319) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78320 && (row * 640 + col) <= 78333) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78334 && (row * 640 + col) <= 78361) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78362 && (row * 640 + col) <= 78375) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78376 && (row * 640 + col) <= 78403) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78404 && (row * 640 + col) <= 78417) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78418 && (row * 640 + col) <= 78424) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78425 && (row * 640 + col) <= 78438) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78439 && (row * 640 + col) <= 78452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78453 && (row * 640 + col) <= 78466) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78467 && (row * 640 + col) <= 78480) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78481 && (row * 640 + col) <= 78494) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78495 && (row * 640 + col) <= 78522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78523 && (row * 640 + col) <= 78536) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78537 && (row * 640 + col) <= 78543) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78544 && (row * 640 + col) <= 78557) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78558 && (row * 640 + col) <= 78564) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78565 && (row * 640 + col) <= 78578) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78579 && (row * 640 + col) <= 78606) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78607 && (row * 640 + col) <= 78620) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78621 && (row * 640 + col) <= 78627) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78628 && (row * 640 + col) <= 78641) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78642 && (row * 640 + col) <= 78682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78683 && (row * 640 + col) <= 78754) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 78755 && (row * 640 + col) <= 78791) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78792 && (row * 640 + col) <= 78805) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78806 && (row * 640 + col) <= 78833) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78834 && (row * 640 + col) <= 78847) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78848 && (row * 640 + col) <= 78854) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78855 && (row * 640 + col) <= 78868) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78869 && (row * 640 + col) <= 78875) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78876 && (row * 640 + col) <= 78889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78890 && (row * 640 + col) <= 78896) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78897 && (row * 640 + col) <= 78910) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78911 && (row * 640 + col) <= 78924) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78925 && (row * 640 + col) <= 78938) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78939 && (row * 640 + col) <= 78959) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78960 && (row * 640 + col) <= 78973) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 78974 && (row * 640 + col) <= 79001) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79002 && (row * 640 + col) <= 79015) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79016 && (row * 640 + col) <= 79043) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79044 && (row * 640 + col) <= 79057) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79058 && (row * 640 + col) <= 79064) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79065 && (row * 640 + col) <= 79078) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79079 && (row * 640 + col) <= 79092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79093 && (row * 640 + col) <= 79106) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79107 && (row * 640 + col) <= 79120) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79121 && (row * 640 + col) <= 79134) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79135 && (row * 640 + col) <= 79162) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79163 && (row * 640 + col) <= 79176) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79177 && (row * 640 + col) <= 79183) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79184 && (row * 640 + col) <= 79197) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79198 && (row * 640 + col) <= 79204) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79205 && (row * 640 + col) <= 79218) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79219 && (row * 640 + col) <= 79246) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79247 && (row * 640 + col) <= 79260) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79261 && (row * 640 + col) <= 79267) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79268 && (row * 640 + col) <= 79281) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79282 && (row * 640 + col) <= 79322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79323 && (row * 640 + col) <= 79394) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 79395 && (row * 640 + col) <= 79431) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79432 && (row * 640 + col) <= 79445) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79446 && (row * 640 + col) <= 79473) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79474 && (row * 640 + col) <= 79487) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79488 && (row * 640 + col) <= 79494) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79495 && (row * 640 + col) <= 79508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79509 && (row * 640 + col) <= 79515) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79516 && (row * 640 + col) <= 79529) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79530 && (row * 640 + col) <= 79536) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79537 && (row * 640 + col) <= 79550) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79551 && (row * 640 + col) <= 79564) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79565 && (row * 640 + col) <= 79578) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79579 && (row * 640 + col) <= 79599) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79600 && (row * 640 + col) <= 79613) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79614 && (row * 640 + col) <= 79641) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79642 && (row * 640 + col) <= 79655) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79656 && (row * 640 + col) <= 79683) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79684 && (row * 640 + col) <= 79697) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79698 && (row * 640 + col) <= 79704) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79705 && (row * 640 + col) <= 79718) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79719 && (row * 640 + col) <= 79732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79733 && (row * 640 + col) <= 79746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79747 && (row * 640 + col) <= 79760) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79761 && (row * 640 + col) <= 79774) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79775 && (row * 640 + col) <= 79802) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79803 && (row * 640 + col) <= 79816) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79817 && (row * 640 + col) <= 79823) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79824 && (row * 640 + col) <= 79837) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79838 && (row * 640 + col) <= 79844) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79845 && (row * 640 + col) <= 79858) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79859 && (row * 640 + col) <= 79886) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79887 && (row * 640 + col) <= 79900) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79901 && (row * 640 + col) <= 79907) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79908 && (row * 640 + col) <= 79921) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 79922 && (row * 640 + col) <= 79962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79963 && (row * 640 + col) <= 80034) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 80035 && (row * 640 + col) <= 80071) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80072 && (row * 640 + col) <= 80085) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80086 && (row * 640 + col) <= 80113) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80114 && (row * 640 + col) <= 80127) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80128 && (row * 640 + col) <= 80134) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80135 && (row * 640 + col) <= 80148) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80149 && (row * 640 + col) <= 80155) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80156 && (row * 640 + col) <= 80169) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80170 && (row * 640 + col) <= 80176) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80177 && (row * 640 + col) <= 80190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80191 && (row * 640 + col) <= 80204) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80205 && (row * 640 + col) <= 80218) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80219 && (row * 640 + col) <= 80239) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80240 && (row * 640 + col) <= 80253) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80254 && (row * 640 + col) <= 80281) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80282 && (row * 640 + col) <= 80295) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80296 && (row * 640 + col) <= 80323) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80324 && (row * 640 + col) <= 80337) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80338 && (row * 640 + col) <= 80344) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80345 && (row * 640 + col) <= 80358) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80359 && (row * 640 + col) <= 80372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80373 && (row * 640 + col) <= 80386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80387 && (row * 640 + col) <= 80400) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80401 && (row * 640 + col) <= 80414) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80415 && (row * 640 + col) <= 80442) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80443 && (row * 640 + col) <= 80456) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80457 && (row * 640 + col) <= 80463) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80464 && (row * 640 + col) <= 80477) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80478 && (row * 640 + col) <= 80484) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80485 && (row * 640 + col) <= 80498) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80499 && (row * 640 + col) <= 80526) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80527 && (row * 640 + col) <= 80540) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80541 && (row * 640 + col) <= 80547) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80548 && (row * 640 + col) <= 80561) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80562 && (row * 640 + col) <= 80602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80603 && (row * 640 + col) <= 80674) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 80675 && (row * 640 + col) <= 80711) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80712 && (row * 640 + col) <= 80725) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80726 && (row * 640 + col) <= 80753) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80754 && (row * 640 + col) <= 80767) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80768 && (row * 640 + col) <= 80774) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80775 && (row * 640 + col) <= 80788) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80789 && (row * 640 + col) <= 80795) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80796 && (row * 640 + col) <= 80809) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80810 && (row * 640 + col) <= 80816) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80817 && (row * 640 + col) <= 80830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80831 && (row * 640 + col) <= 80844) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80845 && (row * 640 + col) <= 80858) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80859 && (row * 640 + col) <= 80879) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80880 && (row * 640 + col) <= 80893) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80894 && (row * 640 + col) <= 80921) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80922 && (row * 640 + col) <= 80935) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80936 && (row * 640 + col) <= 80963) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80964 && (row * 640 + col) <= 80977) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80978 && (row * 640 + col) <= 80984) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80985 && (row * 640 + col) <= 80998) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 80999 && (row * 640 + col) <= 81012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81013 && (row * 640 + col) <= 81026) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81027 && (row * 640 + col) <= 81040) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81041 && (row * 640 + col) <= 81054) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81055 && (row * 640 + col) <= 81082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81083 && (row * 640 + col) <= 81096) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81097 && (row * 640 + col) <= 81103) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81104 && (row * 640 + col) <= 81117) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81118 && (row * 640 + col) <= 81124) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81125 && (row * 640 + col) <= 81138) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81139 && (row * 640 + col) <= 81166) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81167 && (row * 640 + col) <= 81180) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81181 && (row * 640 + col) <= 81187) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81188 && (row * 640 + col) <= 81201) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81202 && (row * 640 + col) <= 81242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81243 && (row * 640 + col) <= 81314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 81315 && (row * 640 + col) <= 81351) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81352 && (row * 640 + col) <= 81365) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81366 && (row * 640 + col) <= 81393) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81394 && (row * 640 + col) <= 81407) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81408 && (row * 640 + col) <= 81414) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81415 && (row * 640 + col) <= 81428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81429 && (row * 640 + col) <= 81435) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81436 && (row * 640 + col) <= 81449) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81450 && (row * 640 + col) <= 81456) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81457 && (row * 640 + col) <= 81470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81471 && (row * 640 + col) <= 81484) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81485 && (row * 640 + col) <= 81498) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81499 && (row * 640 + col) <= 81519) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81520 && (row * 640 + col) <= 81533) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81534 && (row * 640 + col) <= 81561) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81562 && (row * 640 + col) <= 81575) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81576 && (row * 640 + col) <= 81603) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81604 && (row * 640 + col) <= 81617) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81618 && (row * 640 + col) <= 81624) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81625 && (row * 640 + col) <= 81638) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81639 && (row * 640 + col) <= 81652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81653 && (row * 640 + col) <= 81666) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81667 && (row * 640 + col) <= 81680) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81681 && (row * 640 + col) <= 81694) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81695 && (row * 640 + col) <= 81722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81723 && (row * 640 + col) <= 81736) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81737 && (row * 640 + col) <= 81743) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81744 && (row * 640 + col) <= 81757) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81758 && (row * 640 + col) <= 81764) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81765 && (row * 640 + col) <= 81778) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81779 && (row * 640 + col) <= 81806) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81807 && (row * 640 + col) <= 81820) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81821 && (row * 640 + col) <= 81827) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81828 && (row * 640 + col) <= 81841) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 81842 && (row * 640 + col) <= 81882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81883 && (row * 640 + col) <= 81954) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 81955 && (row * 640 + col) <= 81991) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81992 && (row * 640 + col) <= 82005) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82006 && (row * 640 + col) <= 82033) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82034 && (row * 640 + col) <= 82047) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82048 && (row * 640 + col) <= 82054) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82055 && (row * 640 + col) <= 82068) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82069 && (row * 640 + col) <= 82075) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82076 && (row * 640 + col) <= 82089) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82090 && (row * 640 + col) <= 82096) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82097 && (row * 640 + col) <= 82110) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82111 && (row * 640 + col) <= 82124) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82125 && (row * 640 + col) <= 82138) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82139 && (row * 640 + col) <= 82159) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82160 && (row * 640 + col) <= 82173) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82174 && (row * 640 + col) <= 82201) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82202 && (row * 640 + col) <= 82215) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82216 && (row * 640 + col) <= 82243) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82244 && (row * 640 + col) <= 82257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82258 && (row * 640 + col) <= 82264) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82265 && (row * 640 + col) <= 82278) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82279 && (row * 640 + col) <= 82292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82293 && (row * 640 + col) <= 82306) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82307 && (row * 640 + col) <= 82320) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82321 && (row * 640 + col) <= 82334) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82335 && (row * 640 + col) <= 82362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82363 && (row * 640 + col) <= 82376) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82377 && (row * 640 + col) <= 82383) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82384 && (row * 640 + col) <= 82397) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82398 && (row * 640 + col) <= 82404) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82405 && (row * 640 + col) <= 82418) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82419 && (row * 640 + col) <= 82446) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82447 && (row * 640 + col) <= 82460) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82461 && (row * 640 + col) <= 82467) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82468 && (row * 640 + col) <= 82481) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82482 && (row * 640 + col) <= 82522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82523 && (row * 640 + col) <= 82594) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 82595 && (row * 640 + col) <= 82631) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82632 && (row * 640 + col) <= 82645) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82646 && (row * 640 + col) <= 82673) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82674 && (row * 640 + col) <= 82687) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82688 && (row * 640 + col) <= 82694) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82695 && (row * 640 + col) <= 82708) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82709 && (row * 640 + col) <= 82715) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82716 && (row * 640 + col) <= 82729) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82730 && (row * 640 + col) <= 82736) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82737 && (row * 640 + col) <= 82750) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82751 && (row * 640 + col) <= 82764) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82765 && (row * 640 + col) <= 82778) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82779 && (row * 640 + col) <= 82799) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82800 && (row * 640 + col) <= 82813) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82814 && (row * 640 + col) <= 82841) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82842 && (row * 640 + col) <= 82855) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82856 && (row * 640 + col) <= 82883) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82884 && (row * 640 + col) <= 82897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82898 && (row * 640 + col) <= 82904) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82905 && (row * 640 + col) <= 82918) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82919 && (row * 640 + col) <= 82932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82933 && (row * 640 + col) <= 82946) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82947 && (row * 640 + col) <= 82960) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82961 && (row * 640 + col) <= 82974) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 82975 && (row * 640 + col) <= 83002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83003 && (row * 640 + col) <= 83016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83017 && (row * 640 + col) <= 83023) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83024 && (row * 640 + col) <= 83037) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83038 && (row * 640 + col) <= 83044) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83045 && (row * 640 + col) <= 83058) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83059 && (row * 640 + col) <= 83086) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83087 && (row * 640 + col) <= 83100) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83101 && (row * 640 + col) <= 83107) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83108 && (row * 640 + col) <= 83121) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83122 && (row * 640 + col) <= 83162) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83163 && (row * 640 + col) <= 83234) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 83235 && (row * 640 + col) <= 83271) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83272 && (row * 640 + col) <= 83285) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83286 && (row * 640 + col) <= 83313) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83314 && (row * 640 + col) <= 83327) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83328 && (row * 640 + col) <= 83334) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83335 && (row * 640 + col) <= 83348) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83349 && (row * 640 + col) <= 83355) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83356 && (row * 640 + col) <= 83369) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83370 && (row * 640 + col) <= 83376) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83377 && (row * 640 + col) <= 83390) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83391 && (row * 640 + col) <= 83404) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83405 && (row * 640 + col) <= 83418) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83419 && (row * 640 + col) <= 83439) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83440 && (row * 640 + col) <= 83453) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83454 && (row * 640 + col) <= 83481) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83482 && (row * 640 + col) <= 83495) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83496 && (row * 640 + col) <= 83502) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83503 && (row * 640 + col) <= 83516) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83517 && (row * 640 + col) <= 83523) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83524 && (row * 640 + col) <= 83537) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83538 && (row * 640 + col) <= 83544) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83545 && (row * 640 + col) <= 83558) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83559 && (row * 640 + col) <= 83572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83573 && (row * 640 + col) <= 83586) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83587 && (row * 640 + col) <= 83600) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83601 && (row * 640 + col) <= 83614) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83615 && (row * 640 + col) <= 83621) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83622 && (row * 640 + col) <= 83635) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83636 && (row * 640 + col) <= 83642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83643 && (row * 640 + col) <= 83656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83657 && (row * 640 + col) <= 83663) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83664 && (row * 640 + col) <= 83677) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83678 && (row * 640 + col) <= 83684) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83685 && (row * 640 + col) <= 83698) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83699 && (row * 640 + col) <= 83705) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83706 && (row * 640 + col) <= 83719) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83720 && (row * 640 + col) <= 83726) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83727 && (row * 640 + col) <= 83740) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83741 && (row * 640 + col) <= 83747) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83748 && (row * 640 + col) <= 83761) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83762 && (row * 640 + col) <= 83802) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83803 && (row * 640 + col) <= 83874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 83875 && (row * 640 + col) <= 83911) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83912 && (row * 640 + col) <= 83925) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83926 && (row * 640 + col) <= 83953) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83954 && (row * 640 + col) <= 83967) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83968 && (row * 640 + col) <= 83974) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83975 && (row * 640 + col) <= 83988) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 83989 && (row * 640 + col) <= 83995) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83996 && (row * 640 + col) <= 84009) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84010 && (row * 640 + col) <= 84016) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84017 && (row * 640 + col) <= 84030) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84031 && (row * 640 + col) <= 84044) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84045 && (row * 640 + col) <= 84058) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84059 && (row * 640 + col) <= 84079) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84080 && (row * 640 + col) <= 84093) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84094 && (row * 640 + col) <= 84121) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84122 && (row * 640 + col) <= 84135) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84136 && (row * 640 + col) <= 84142) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84143 && (row * 640 + col) <= 84156) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84157 && (row * 640 + col) <= 84163) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84164 && (row * 640 + col) <= 84177) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84178 && (row * 640 + col) <= 84184) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84185 && (row * 640 + col) <= 84198) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84199 && (row * 640 + col) <= 84212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84213 && (row * 640 + col) <= 84226) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84227 && (row * 640 + col) <= 84240) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84241 && (row * 640 + col) <= 84254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84255 && (row * 640 + col) <= 84261) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84262 && (row * 640 + col) <= 84275) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84276 && (row * 640 + col) <= 84282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84283 && (row * 640 + col) <= 84296) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84297 && (row * 640 + col) <= 84303) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84304 && (row * 640 + col) <= 84317) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84318 && (row * 640 + col) <= 84324) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84325 && (row * 640 + col) <= 84338) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84339 && (row * 640 + col) <= 84345) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84346 && (row * 640 + col) <= 84359) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84360 && (row * 640 + col) <= 84366) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84367 && (row * 640 + col) <= 84380) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84381 && (row * 640 + col) <= 84387) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84388 && (row * 640 + col) <= 84401) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84402 && (row * 640 + col) <= 84442) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84443 && (row * 640 + col) <= 84514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 84515 && (row * 640 + col) <= 84551) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84552 && (row * 640 + col) <= 84565) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84566 && (row * 640 + col) <= 84593) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84594 && (row * 640 + col) <= 84607) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84608 && (row * 640 + col) <= 84614) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84615 && (row * 640 + col) <= 84628) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84629 && (row * 640 + col) <= 84635) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84636 && (row * 640 + col) <= 84649) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84650 && (row * 640 + col) <= 84656) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84657 && (row * 640 + col) <= 84670) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84671 && (row * 640 + col) <= 84684) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84685 && (row * 640 + col) <= 84698) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84699 && (row * 640 + col) <= 84719) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84720 && (row * 640 + col) <= 84733) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84734 && (row * 640 + col) <= 84761) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84762 && (row * 640 + col) <= 84775) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84776 && (row * 640 + col) <= 84782) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84783 && (row * 640 + col) <= 84796) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84797 && (row * 640 + col) <= 84803) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84804 && (row * 640 + col) <= 84817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84818 && (row * 640 + col) <= 84824) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84825 && (row * 640 + col) <= 84838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84839 && (row * 640 + col) <= 84852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84853 && (row * 640 + col) <= 84866) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84867 && (row * 640 + col) <= 84880) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84881 && (row * 640 + col) <= 84894) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84895 && (row * 640 + col) <= 84901) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84902 && (row * 640 + col) <= 84915) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84916 && (row * 640 + col) <= 84922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84923 && (row * 640 + col) <= 84936) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84937 && (row * 640 + col) <= 84943) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84944 && (row * 640 + col) <= 84957) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84958 && (row * 640 + col) <= 84964) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84965 && (row * 640 + col) <= 84978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 84979 && (row * 640 + col) <= 84985) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84986 && (row * 640 + col) <= 84999) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85000 && (row * 640 + col) <= 85006) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85007 && (row * 640 + col) <= 85020) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85021 && (row * 640 + col) <= 85027) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85028 && (row * 640 + col) <= 85041) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85042 && (row * 640 + col) <= 85082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85083 && (row * 640 + col) <= 85154) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 85155 && (row * 640 + col) <= 85191) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85192 && (row * 640 + col) <= 85205) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85206 && (row * 640 + col) <= 85233) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85234 && (row * 640 + col) <= 85247) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85248 && (row * 640 + col) <= 85254) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85255 && (row * 640 + col) <= 85268) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85269 && (row * 640 + col) <= 85275) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85276 && (row * 640 + col) <= 85289) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85290 && (row * 640 + col) <= 85296) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85297 && (row * 640 + col) <= 85310) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85311 && (row * 640 + col) <= 85324) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85325 && (row * 640 + col) <= 85338) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85339 && (row * 640 + col) <= 85359) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85360 && (row * 640 + col) <= 85373) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85374 && (row * 640 + col) <= 85401) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85402 && (row * 640 + col) <= 85415) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85416 && (row * 640 + col) <= 85422) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85423 && (row * 640 + col) <= 85436) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85437 && (row * 640 + col) <= 85443) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85444 && (row * 640 + col) <= 85457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85458 && (row * 640 + col) <= 85464) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85465 && (row * 640 + col) <= 85478) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85479 && (row * 640 + col) <= 85492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85493 && (row * 640 + col) <= 85506) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85507 && (row * 640 + col) <= 85520) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85521 && (row * 640 + col) <= 85534) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85535 && (row * 640 + col) <= 85541) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85542 && (row * 640 + col) <= 85555) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85556 && (row * 640 + col) <= 85562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85563 && (row * 640 + col) <= 85576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85577 && (row * 640 + col) <= 85583) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85584 && (row * 640 + col) <= 85597) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85598 && (row * 640 + col) <= 85604) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85605 && (row * 640 + col) <= 85618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85619 && (row * 640 + col) <= 85625) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85626 && (row * 640 + col) <= 85639) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85640 && (row * 640 + col) <= 85646) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85647 && (row * 640 + col) <= 85660) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85661 && (row * 640 + col) <= 85667) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85668 && (row * 640 + col) <= 85681) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85682 && (row * 640 + col) <= 85722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85723 && (row * 640 + col) <= 85794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 85795 && (row * 640 + col) <= 85831) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85832 && (row * 640 + col) <= 85845) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85846 && (row * 640 + col) <= 85873) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85874 && (row * 640 + col) <= 85887) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85888 && (row * 640 + col) <= 85894) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85895 && (row * 640 + col) <= 85908) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85909 && (row * 640 + col) <= 85915) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85916 && (row * 640 + col) <= 85929) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85930 && (row * 640 + col) <= 85936) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85937 && (row * 640 + col) <= 85950) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85951 && (row * 640 + col) <= 85964) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85965 && (row * 640 + col) <= 85978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 85979 && (row * 640 + col) <= 85999) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86000 && (row * 640 + col) <= 86013) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86014 && (row * 640 + col) <= 86041) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86042 && (row * 640 + col) <= 86055) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86056 && (row * 640 + col) <= 86062) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86063 && (row * 640 + col) <= 86076) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86077 && (row * 640 + col) <= 86083) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86084 && (row * 640 + col) <= 86097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86098 && (row * 640 + col) <= 86104) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86105 && (row * 640 + col) <= 86118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86119 && (row * 640 + col) <= 86132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86133 && (row * 640 + col) <= 86146) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86147 && (row * 640 + col) <= 86160) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86161 && (row * 640 + col) <= 86174) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86175 && (row * 640 + col) <= 86181) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86182 && (row * 640 + col) <= 86195) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86196 && (row * 640 + col) <= 86202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86203 && (row * 640 + col) <= 86216) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86217 && (row * 640 + col) <= 86223) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86224 && (row * 640 + col) <= 86237) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86238 && (row * 640 + col) <= 86244) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86245 && (row * 640 + col) <= 86258) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86259 && (row * 640 + col) <= 86265) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86266 && (row * 640 + col) <= 86279) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86280 && (row * 640 + col) <= 86286) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86287 && (row * 640 + col) <= 86300) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86301 && (row * 640 + col) <= 86307) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86308 && (row * 640 + col) <= 86321) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86322 && (row * 640 + col) <= 86362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86363 && (row * 640 + col) <= 86434) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 86435 && (row * 640 + col) <= 86471) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86472 && (row * 640 + col) <= 86485) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86486 && (row * 640 + col) <= 86513) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86514 && (row * 640 + col) <= 86527) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86528 && (row * 640 + col) <= 86534) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86535 && (row * 640 + col) <= 86548) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86549 && (row * 640 + col) <= 86555) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86556 && (row * 640 + col) <= 86569) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86570 && (row * 640 + col) <= 86576) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86577 && (row * 640 + col) <= 86590) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86591 && (row * 640 + col) <= 86604) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86605 && (row * 640 + col) <= 86618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86619 && (row * 640 + col) <= 86639) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86640 && (row * 640 + col) <= 86653) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86654 && (row * 640 + col) <= 86681) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86682 && (row * 640 + col) <= 86695) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86696 && (row * 640 + col) <= 86702) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86703 && (row * 640 + col) <= 86716) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86717 && (row * 640 + col) <= 86723) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86724 && (row * 640 + col) <= 86737) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86738 && (row * 640 + col) <= 86744) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86745 && (row * 640 + col) <= 86758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86759 && (row * 640 + col) <= 86772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86773 && (row * 640 + col) <= 86786) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86787 && (row * 640 + col) <= 86800) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86801 && (row * 640 + col) <= 86814) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86815 && (row * 640 + col) <= 86821) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86822 && (row * 640 + col) <= 86835) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86836 && (row * 640 + col) <= 86842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86843 && (row * 640 + col) <= 86856) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86857 && (row * 640 + col) <= 86863) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86864 && (row * 640 + col) <= 86877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86878 && (row * 640 + col) <= 86884) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86885 && (row * 640 + col) <= 86898) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86899 && (row * 640 + col) <= 86905) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86906 && (row * 640 + col) <= 86919) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86920 && (row * 640 + col) <= 86926) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86927 && (row * 640 + col) <= 86940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86941 && (row * 640 + col) <= 86947) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86948 && (row * 640 + col) <= 86961) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 86962 && (row * 640 + col) <= 87002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87003 && (row * 640 + col) <= 87074) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87075 && (row * 640 + col) <= 87111) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87112 && (row * 640 + col) <= 87125) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87126 && (row * 640 + col) <= 87153) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87154 && (row * 640 + col) <= 87167) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87168 && (row * 640 + col) <= 87174) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87175 && (row * 640 + col) <= 87188) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87189 && (row * 640 + col) <= 87195) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87196 && (row * 640 + col) <= 87209) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87210 && (row * 640 + col) <= 87216) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87217 && (row * 640 + col) <= 87230) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87231 && (row * 640 + col) <= 87244) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87245 && (row * 640 + col) <= 87258) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87259 && (row * 640 + col) <= 87279) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87280 && (row * 640 + col) <= 87293) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87294 && (row * 640 + col) <= 87321) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87322 && (row * 640 + col) <= 87335) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87336 && (row * 640 + col) <= 87342) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87343 && (row * 640 + col) <= 87356) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87357 && (row * 640 + col) <= 87363) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87364 && (row * 640 + col) <= 87377) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87378 && (row * 640 + col) <= 87384) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87385 && (row * 640 + col) <= 87398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87399 && (row * 640 + col) <= 87412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87413 && (row * 640 + col) <= 87426) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87427 && (row * 640 + col) <= 87440) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87441 && (row * 640 + col) <= 87454) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87455 && (row * 640 + col) <= 87461) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87462 && (row * 640 + col) <= 87475) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87476 && (row * 640 + col) <= 87482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87483 && (row * 640 + col) <= 87496) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87497 && (row * 640 + col) <= 87503) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87504 && (row * 640 + col) <= 87517) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87518 && (row * 640 + col) <= 87524) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87525 && (row * 640 + col) <= 87538) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87539 && (row * 640 + col) <= 87545) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87546 && (row * 640 + col) <= 87559) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87560 && (row * 640 + col) <= 87566) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87567 && (row * 640 + col) <= 87580) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87581 && (row * 640 + col) <= 87587) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87588 && (row * 640 + col) <= 87601) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87602 && (row * 640 + col) <= 87642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87643 && (row * 640 + col) <= 87714) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87715 && (row * 640 + col) <= 87751) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87752 && (row * 640 + col) <= 87765) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87766 && (row * 640 + col) <= 87793) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87794 && (row * 640 + col) <= 87807) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87808 && (row * 640 + col) <= 87814) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87815 && (row * 640 + col) <= 87828) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87829 && (row * 640 + col) <= 87835) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87836 && (row * 640 + col) <= 87870) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87871 && (row * 640 + col) <= 87877) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87878 && (row * 640 + col) <= 87905) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87906 && (row * 640 + col) <= 87919) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87920 && (row * 640 + col) <= 87933) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87934 && (row * 640 + col) <= 87961) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87962 && (row * 640 + col) <= 87996) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 87997 && (row * 640 + col) <= 88003) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88004 && (row * 640 + col) <= 88017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88018 && (row * 640 + col) <= 88024) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88025 && (row * 640 + col) <= 88038) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88039 && (row * 640 + col) <= 88052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88053 && (row * 640 + col) <= 88066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88067 && (row * 640 + col) <= 88080) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88081 && (row * 640 + col) <= 88115) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88116 && (row * 640 + col) <= 88122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88123 && (row * 640 + col) <= 88136) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88137 && (row * 640 + col) <= 88143) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88144 && (row * 640 + col) <= 88157) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88158 && (row * 640 + col) <= 88164) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88165 && (row * 640 + col) <= 88199) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88200 && (row * 640 + col) <= 88206) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88207 && (row * 640 + col) <= 88220) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88221 && (row * 640 + col) <= 88227) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88228 && (row * 640 + col) <= 88241) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88242 && (row * 640 + col) <= 88282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88283 && (row * 640 + col) <= 88354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88355 && (row * 640 + col) <= 88391) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88392 && (row * 640 + col) <= 88405) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88406 && (row * 640 + col) <= 88433) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88434 && (row * 640 + col) <= 88447) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88448 && (row * 640 + col) <= 88454) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88455 && (row * 640 + col) <= 88468) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88469 && (row * 640 + col) <= 88475) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88476 && (row * 640 + col) <= 88510) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88511 && (row * 640 + col) <= 88517) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88518 && (row * 640 + col) <= 88545) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88546 && (row * 640 + col) <= 88559) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88560 && (row * 640 + col) <= 88573) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88574 && (row * 640 + col) <= 88601) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88602 && (row * 640 + col) <= 88636) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88637 && (row * 640 + col) <= 88643) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88644 && (row * 640 + col) <= 88657) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88658 && (row * 640 + col) <= 88664) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88665 && (row * 640 + col) <= 88678) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88679 && (row * 640 + col) <= 88692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88693 && (row * 640 + col) <= 88706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88707 && (row * 640 + col) <= 88720) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88721 && (row * 640 + col) <= 88755) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88756 && (row * 640 + col) <= 88762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88763 && (row * 640 + col) <= 88776) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88777 && (row * 640 + col) <= 88783) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88784 && (row * 640 + col) <= 88797) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88798 && (row * 640 + col) <= 88804) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88805 && (row * 640 + col) <= 88839) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88840 && (row * 640 + col) <= 88846) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88847 && (row * 640 + col) <= 88860) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88861 && (row * 640 + col) <= 88867) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88868 && (row * 640 + col) <= 88881) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 88882 && (row * 640 + col) <= 88922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88923 && (row * 640 + col) <= 88994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88995 && (row * 640 + col) <= 89031) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89032 && (row * 640 + col) <= 89045) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89046 && (row * 640 + col) <= 89073) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89074 && (row * 640 + col) <= 89087) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89088 && (row * 640 + col) <= 89094) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89095 && (row * 640 + col) <= 89108) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89109 && (row * 640 + col) <= 89115) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89116 && (row * 640 + col) <= 89150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89151 && (row * 640 + col) <= 89157) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89158 && (row * 640 + col) <= 89185) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89186 && (row * 640 + col) <= 89199) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89200 && (row * 640 + col) <= 89213) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89214 && (row * 640 + col) <= 89241) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89242 && (row * 640 + col) <= 89276) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89277 && (row * 640 + col) <= 89283) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89284 && (row * 640 + col) <= 89297) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89298 && (row * 640 + col) <= 89304) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89305 && (row * 640 + col) <= 89318) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89319 && (row * 640 + col) <= 89332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89333 && (row * 640 + col) <= 89346) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89347 && (row * 640 + col) <= 89360) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89361 && (row * 640 + col) <= 89395) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89396 && (row * 640 + col) <= 89402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89403 && (row * 640 + col) <= 89416) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89417 && (row * 640 + col) <= 89423) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89424 && (row * 640 + col) <= 89437) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89438 && (row * 640 + col) <= 89444) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89445 && (row * 640 + col) <= 89479) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89480 && (row * 640 + col) <= 89486) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89487 && (row * 640 + col) <= 89500) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89501 && (row * 640 + col) <= 89507) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89508 && (row * 640 + col) <= 89521) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89522 && (row * 640 + col) <= 89562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89563 && (row * 640 + col) <= 89634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 89635 && (row * 640 + col) <= 89671) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89672 && (row * 640 + col) <= 89685) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89686 && (row * 640 + col) <= 89713) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89714 && (row * 640 + col) <= 89727) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89728 && (row * 640 + col) <= 89734) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89735 && (row * 640 + col) <= 89748) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89749 && (row * 640 + col) <= 89755) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89756 && (row * 640 + col) <= 89790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89791 && (row * 640 + col) <= 89797) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89798 && (row * 640 + col) <= 89825) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89826 && (row * 640 + col) <= 89839) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89840 && (row * 640 + col) <= 89853) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89854 && (row * 640 + col) <= 89881) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89882 && (row * 640 + col) <= 89916) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89917 && (row * 640 + col) <= 89923) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89924 && (row * 640 + col) <= 89937) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89938 && (row * 640 + col) <= 89944) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89945 && (row * 640 + col) <= 89958) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89959 && (row * 640 + col) <= 89972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89973 && (row * 640 + col) <= 89986) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 89987 && (row * 640 + col) <= 90000) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90001 && (row * 640 + col) <= 90035) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90036 && (row * 640 + col) <= 90042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90043 && (row * 640 + col) <= 90056) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90057 && (row * 640 + col) <= 90063) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90064 && (row * 640 + col) <= 90077) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90078 && (row * 640 + col) <= 90084) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90085 && (row * 640 + col) <= 90119) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90120 && (row * 640 + col) <= 90126) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90127 && (row * 640 + col) <= 90140) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90141 && (row * 640 + col) <= 90147) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90148 && (row * 640 + col) <= 90161) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90162 && (row * 640 + col) <= 90202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90203 && (row * 640 + col) <= 90274) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 90275 && (row * 640 + col) <= 90311) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90312 && (row * 640 + col) <= 90325) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90326 && (row * 640 + col) <= 90353) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90354 && (row * 640 + col) <= 90367) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90368 && (row * 640 + col) <= 90374) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90375 && (row * 640 + col) <= 90388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90389 && (row * 640 + col) <= 90395) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90396 && (row * 640 + col) <= 90430) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90431 && (row * 640 + col) <= 90437) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90438 && (row * 640 + col) <= 90465) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90466 && (row * 640 + col) <= 90479) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90480 && (row * 640 + col) <= 90493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90494 && (row * 640 + col) <= 90521) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90522 && (row * 640 + col) <= 90556) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90557 && (row * 640 + col) <= 90563) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90564 && (row * 640 + col) <= 90577) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90578 && (row * 640 + col) <= 90584) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90585 && (row * 640 + col) <= 90598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90599 && (row * 640 + col) <= 90612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90613 && (row * 640 + col) <= 90626) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90627 && (row * 640 + col) <= 90640) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90641 && (row * 640 + col) <= 90675) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90676 && (row * 640 + col) <= 90682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90683 && (row * 640 + col) <= 90696) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90697 && (row * 640 + col) <= 90703) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90704 && (row * 640 + col) <= 90717) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90718 && (row * 640 + col) <= 90724) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90725 && (row * 640 + col) <= 90759) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90760 && (row * 640 + col) <= 90766) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90767 && (row * 640 + col) <= 90780) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90781 && (row * 640 + col) <= 90787) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90788 && (row * 640 + col) <= 90801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90802 && (row * 640 + col) <= 90842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90843 && (row * 640 + col) <= 90914) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 90915 && (row * 640 + col) <= 90951) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90952 && (row * 640 + col) <= 90965) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 90966 && (row * 640 + col) <= 90993) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90994 && (row * 640 + col) <= 91007) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91008 && (row * 640 + col) <= 91014) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91015 && (row * 640 + col) <= 91028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91029 && (row * 640 + col) <= 91035) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91036 && (row * 640 + col) <= 91070) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91071 && (row * 640 + col) <= 91077) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91078 && (row * 640 + col) <= 91105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91106 && (row * 640 + col) <= 91119) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91120 && (row * 640 + col) <= 91133) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91134 && (row * 640 + col) <= 91161) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91162 && (row * 640 + col) <= 91196) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91197 && (row * 640 + col) <= 91203) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91204 && (row * 640 + col) <= 91217) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91218 && (row * 640 + col) <= 91224) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91225 && (row * 640 + col) <= 91238) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91239 && (row * 640 + col) <= 91252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91253 && (row * 640 + col) <= 91266) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91267 && (row * 640 + col) <= 91280) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91281 && (row * 640 + col) <= 91315) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91316 && (row * 640 + col) <= 91322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91323 && (row * 640 + col) <= 91336) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91337 && (row * 640 + col) <= 91343) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91344 && (row * 640 + col) <= 91357) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91358 && (row * 640 + col) <= 91364) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91365 && (row * 640 + col) <= 91399) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91400 && (row * 640 + col) <= 91406) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91407 && (row * 640 + col) <= 91420) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91421 && (row * 640 + col) <= 91427) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91428 && (row * 640 + col) <= 91441) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91442 && (row * 640 + col) <= 91482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91483 && (row * 640 + col) <= 91554) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 91555 && (row * 640 + col) <= 91591) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91592 && (row * 640 + col) <= 91605) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91606 && (row * 640 + col) <= 91633) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91634 && (row * 640 + col) <= 91647) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91648 && (row * 640 + col) <= 91654) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91655 && (row * 640 + col) <= 91668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91669 && (row * 640 + col) <= 91675) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91676 && (row * 640 + col) <= 91710) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91711 && (row * 640 + col) <= 91717) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91718 && (row * 640 + col) <= 91745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91746 && (row * 640 + col) <= 91759) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91760 && (row * 640 + col) <= 91773) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91774 && (row * 640 + col) <= 91801) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91802 && (row * 640 + col) <= 91836) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91837 && (row * 640 + col) <= 91843) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91844 && (row * 640 + col) <= 91857) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91858 && (row * 640 + col) <= 91864) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91865 && (row * 640 + col) <= 91878) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91879 && (row * 640 + col) <= 91892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91893 && (row * 640 + col) <= 91906) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91907 && (row * 640 + col) <= 91920) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91921 && (row * 640 + col) <= 91955) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91956 && (row * 640 + col) <= 91962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91963 && (row * 640 + col) <= 91976) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91977 && (row * 640 + col) <= 91983) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91984 && (row * 640 + col) <= 91997) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 91998 && (row * 640 + col) <= 92004) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 92005 && (row * 640 + col) <= 92039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92040 && (row * 640 + col) <= 92046) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 92047 && (row * 640 + col) <= 92060) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92061 && (row * 640 + col) <= 92067) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 92068 && (row * 640 + col) <= 92081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 92082 && (row * 640 + col) <= 92122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 92123 && (row * 640 + col) <= 92194) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 92195 && (row * 640 + col) <= 92762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 92763 && (row * 640 + col) <= 92834) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 92835 && (row * 640 + col) <= 93402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 93403 && (row * 640 + col) <= 93474) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 93475 && (row * 640 + col) <= 94042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 94043 && (row * 640 + col) <= 94114) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 94115 && (row * 640 + col) <= 94682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 94683 && (row * 640 + col) <= 94754) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 94755 && (row * 640 + col) <= 95322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 95323 && (row * 640 + col) <= 95394) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 95395 && (row * 640 + col) <= 95962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 95963 && (row * 640 + col) <= 96034) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96035 && (row * 640 + col) <= 96602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 96603 && (row * 640 + col) <= 96674) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96675 && (row * 640 + col) <= 97242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97243 && (row * 640 + col) <= 97314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97315 && (row * 640 + col) <= 97882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97883 && (row * 640 + col) <= 97954) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97955 && (row * 640 + col) <= 98522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98523 && (row * 640 + col) <= 98594) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98595 && (row * 640 + col) <= 99162) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99163 && (row * 640 + col) <= 99234) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99235 && (row * 640 + col) <= 99802) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99803 && (row * 640 + col) <= 99874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99875 && (row * 640 + col) <= 100442) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100443 && (row * 640 + col) <= 100514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100515 && (row * 640 + col) <= 101082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101083 && (row * 640 + col) <= 101154) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101155 && (row * 640 + col) <= 101722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101723 && (row * 640 + col) <= 101794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101795 && (row * 640 + col) <= 102362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102363 && (row * 640 + col) <= 102434) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102435 && (row * 640 + col) <= 103002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103003 && (row * 640 + col) <= 103074) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103075 && (row * 640 + col) <= 103642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103643 && (row * 640 + col) <= 103714) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103715 && (row * 640 + col) <= 104282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104283 && (row * 640 + col) <= 104354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104355 && (row * 640 + col) <= 104922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104923 && (row * 640 + col) <= 104994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104995 && (row * 640 + col) <= 105562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105563 && (row * 640 + col) <= 105634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105635 && (row * 640 + col) <= 106202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106203 && (row * 640 + col) <= 106274) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106275 && (row * 640 + col) <= 106842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106843 && (row * 640 + col) <= 106914) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106915 && (row * 640 + col) <= 107482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107483 && (row * 640 + col) <= 107554) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107555 && (row * 640 + col) <= 108122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108123 && (row * 640 + col) <= 108194) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108195 && (row * 640 + col) <= 108762) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108763 && (row * 640 + col) <= 108834) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108835 && (row * 640 + col) <= 109402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109403 && (row * 640 + col) <= 109474) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109475 && (row * 640 + col) <= 110042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110043 && (row * 640 + col) <= 110114) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110115 && (row * 640 + col) <= 110682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110683 && (row * 640 + col) <= 110754) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110755 && (row * 640 + col) <= 111322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111323 && (row * 640 + col) <= 111394) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111395 && (row * 640 + col) <= 111396) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111397 && (row * 640 + col) <= 111400) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 111401 && (row * 640 + col) <= 111956) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111957 && (row * 640 + col) <= 111958) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 111959 && (row * 640 + col) <= 111962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111963 && (row * 640 + col) <= 112034) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112035 && (row * 640 + col) <= 112035) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112036 && (row * 640 + col) <= 112036) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 112037 && (row * 640 + col) <= 112040) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 112041 && (row * 640 + col) <= 112041) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 112042 && (row * 640 + col) <= 112595) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112596 && (row * 640 + col) <= 112596) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 112597 && (row * 640 + col) <= 112598) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 112599 && (row * 640 + col) <= 112599) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 112600 && (row * 640 + col) <= 112602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112603 && (row * 640 + col) <= 112674) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112675 && (row * 640 + col) <= 112675) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112676 && (row * 640 + col) <= 112676) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 112677 && (row * 640 + col) <= 112680) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 112681 && (row * 640 + col) <= 112681) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 112682 && (row * 640 + col) <= 113235) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113236 && (row * 640 + col) <= 113236) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113237 && (row * 640 + col) <= 113239) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 113240 && (row * 640 + col) <= 113240) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113241 && (row * 640 + col) <= 113242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113243 && (row * 640 + col) <= 113310) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113311 && (row * 640 + col) <= 113312) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113313 && (row * 640 + col) <= 113314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113315 && (row * 640 + col) <= 113316) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113317 && (row * 640 + col) <= 113320) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 113321 && (row * 640 + col) <= 113322) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113323 && (row * 640 + col) <= 113324) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113325 && (row * 640 + col) <= 113326) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113327 && (row * 640 + col) <= 113875) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113876 && (row * 640 + col) <= 113876) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113877 && (row * 640 + col) <= 113879) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 113880 && (row * 640 + col) <= 113880) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113881 && (row * 640 + col) <= 113882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113883 && (row * 640 + col) <= 113883) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113884 && (row * 640 + col) <= 113886) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113887 && (row * 640 + col) <= 113949) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113950 && (row * 640 + col) <= 113950) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113951 && (row * 640 + col) <= 113952) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 113953 && (row * 640 + col) <= 113953) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113954 && (row * 640 + col) <= 113954) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113955 && (row * 640 + col) <= 113955) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113956 && (row * 640 + col) <= 113961) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 113962 && (row * 640 + col) <= 113962) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113963 && (row * 640 + col) <= 113963) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113964 && (row * 640 + col) <= 113964) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113965 && (row * 640 + col) <= 113966) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 113967 && (row * 640 + col) <= 113967) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 113968 && (row * 640 + col) <= 114509) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114510 && (row * 640 + col) <= 114512) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114513 && (row * 640 + col) <= 114515) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114516 && (row * 640 + col) <= 114516) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114517 && (row * 640 + col) <= 114519) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 114520 && (row * 640 + col) <= 114520) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114521 && (row * 640 + col) <= 114522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114523 && (row * 640 + col) <= 114523) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114524 && (row * 640 + col) <= 114524) color_data <= 12'b010010110000; else
        if ((row * 640 + col) >= 114525 && (row * 640 + col) <= 114526) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 114527 && (row * 640 + col) <= 114527) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114528 && (row * 640 + col) <= 114589) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114590 && (row * 640 + col) <= 114590) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114591 && (row * 640 + col) <= 114593) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 114594 && (row * 640 + col) <= 114595) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114596 && (row * 640 + col) <= 114601) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 114602 && (row * 640 + col) <= 114603) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114604 && (row * 640 + col) <= 114606) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 114607 && (row * 640 + col) <= 114607) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 114608 && (row * 640 + col) <= 115148) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115149 && (row * 640 + col) <= 115149) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115150 && (row * 640 + col) <= 115152) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 115153 && (row * 640 + col) <= 115154) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115155 && (row * 640 + col) <= 115156) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115157 && (row * 640 + col) <= 115157) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115158 && (row * 640 + col) <= 115159) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 115160 && (row * 640 + col) <= 115160) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115161 && (row * 640 + col) <= 115161) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115162 && (row * 640 + col) <= 115162) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115163 && (row * 640 + col) <= 115165) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 115166 && (row * 640 + col) <= 115166) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115167 && (row * 640 + col) <= 115229) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115230 && (row * 640 + col) <= 115230) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115231 && (row * 640 + col) <= 115234) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 115235 && (row * 640 + col) <= 115235) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115236 && (row * 640 + col) <= 115241) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 115242 && (row * 640 + col) <= 115242) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115243 && (row * 640 + col) <= 115246) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 115247 && (row * 640 + col) <= 115247) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115248 && (row * 640 + col) <= 115788) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115789 && (row * 640 + col) <= 115789) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115790 && (row * 640 + col) <= 115790) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 115791 && (row * 640 + col) <= 115791) color_data <= 12'b010010110000; else
        if ((row * 640 + col) >= 115792 && (row * 640 + col) <= 115794) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 115795 && (row * 640 + col) <= 115795) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115796 && (row * 640 + col) <= 115796) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115797 && (row * 640 + col) <= 115797) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115798 && (row * 640 + col) <= 115799) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 115800 && (row * 640 + col) <= 115801) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115802 && (row * 640 + col) <= 115805) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 115806 && (row * 640 + col) <= 115806) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115807 && (row * 640 + col) <= 115869) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115870 && (row * 640 + col) <= 115870) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115871 && (row * 640 + col) <= 115874) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 115875 && (row * 640 + col) <= 115875) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115876 && (row * 640 + col) <= 115881) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 115882 && (row * 640 + col) <= 115882) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115883 && (row * 640 + col) <= 115886) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 115887 && (row * 640 + col) <= 115887) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 115888 && (row * 640 + col) <= 116429) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116430 && (row * 640 + col) <= 116430) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116431 && (row * 640 + col) <= 116431) color_data <= 12'b010110110001; else
        if ((row * 640 + col) >= 116432 && (row * 640 + col) <= 116435) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 116436 && (row * 640 + col) <= 116437) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116438 && (row * 640 + col) <= 116439) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 116440 && (row * 640 + col) <= 116440) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116441 && (row * 640 + col) <= 116444) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 116445 && (row * 640 + col) <= 116445) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116446 && (row * 640 + col) <= 116510) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116511 && (row * 640 + col) <= 116511) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116512 && (row * 640 + col) <= 116514) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 116515 && (row * 640 + col) <= 116515) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116516 && (row * 640 + col) <= 116521) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 116522 && (row * 640 + col) <= 116522) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116523 && (row * 640 + col) <= 116525) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 116526 && (row * 640 + col) <= 116526) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 116527 && (row * 640 + col) <= 117070) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117071 && (row * 640 + col) <= 117071) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117072 && (row * 640 + col) <= 117072) color_data <= 12'b010110110010; else
        if ((row * 640 + col) >= 117073 && (row * 640 + col) <= 117076) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 117077 && (row * 640 + col) <= 117077) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117078 && (row * 640 + col) <= 117079) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 117080 && (row * 640 + col) <= 117080) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117081 && (row * 640 + col) <= 117084) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 117085 && (row * 640 + col) <= 117085) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117086 && (row * 640 + col) <= 117087) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117088 && (row * 640 + col) <= 117089) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117090 && (row * 640 + col) <= 117146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117147 && (row * 640 + col) <= 117149) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117150 && (row * 640 + col) <= 117150) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117151 && (row * 640 + col) <= 117151) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117152 && (row * 640 + col) <= 117154) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117155 && (row * 640 + col) <= 117155) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117156 && (row * 640 + col) <= 117161) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117162 && (row * 640 + col) <= 117162) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117163 && (row * 640 + col) <= 117165) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117166 && (row * 640 + col) <= 117166) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117167 && (row * 640 + col) <= 117167) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117168 && (row * 640 + col) <= 117171) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117172 && (row * 640 + col) <= 117711) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117712 && (row * 640 + col) <= 117714) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117715 && (row * 640 + col) <= 117716) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 117717 && (row * 640 + col) <= 117717) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117718 && (row * 640 + col) <= 117719) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 117720 && (row * 640 + col) <= 117720) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117721 && (row * 640 + col) <= 117722) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 117723 && (row * 640 + col) <= 117727) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117728 && (row * 640 + col) <= 117728) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 117729 && (row * 640 + col) <= 117729) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117730 && (row * 640 + col) <= 117785) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117786 && (row * 640 + col) <= 117786) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117787 && (row * 640 + col) <= 117789) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117790 && (row * 640 + col) <= 117791) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117792 && (row * 640 + col) <= 117794) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117795 && (row * 640 + col) <= 117796) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117797 && (row * 640 + col) <= 117800) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117801 && (row * 640 + col) <= 117802) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117803 && (row * 640 + col) <= 117804) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117805 && (row * 640 + col) <= 117807) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117808 && (row * 640 + col) <= 117811) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 117812 && (row * 640 + col) <= 117812) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 117813 && (row * 640 + col) <= 118349) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118350 && (row * 640 + col) <= 118351) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118352 && (row * 640 + col) <= 118357) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 118358 && (row * 640 + col) <= 118359) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118360 && (row * 640 + col) <= 118368) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 118369 && (row * 640 + col) <= 118369) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118370 && (row * 640 + col) <= 118424) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118425 && (row * 640 + col) <= 118425) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118426 && (row * 640 + col) <= 118431) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 118432 && (row * 640 + col) <= 118432) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118433 && (row * 640 + col) <= 118435) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 118436 && (row * 640 + col) <= 118436) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118437 && (row * 640 + col) <= 118440) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 118441 && (row * 640 + col) <= 118441) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118442 && (row * 640 + col) <= 118443) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 118444 && (row * 640 + col) <= 118445) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118446 && (row * 640 + col) <= 118450) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 118451 && (row * 640 + col) <= 118451) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118452 && (row * 640 + col) <= 118987) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118988 && (row * 640 + col) <= 118989) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 118990 && (row * 640 + col) <= 119001) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 119002 && (row * 640 + col) <= 119002) color_data <= 12'b000101100000; else
        if ((row * 640 + col) >= 119003 && (row * 640 + col) <= 119006) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 119007 && (row * 640 + col) <= 119008) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119009 && (row * 640 + col) <= 119064) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119065 && (row * 640 + col) <= 119069) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119070 && (row * 640 + col) <= 119072) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119073 && (row * 640 + col) <= 119073) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119074 && (row * 640 + col) <= 119075) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119076 && (row * 640 + col) <= 119077) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119078 && (row * 640 + col) <= 119079) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119080 && (row * 640 + col) <= 119080) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119081 && (row * 640 + col) <= 119082) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119083 && (row * 640 + col) <= 119084) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119085 && (row * 640 + col) <= 119088) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119089 && (row * 640 + col) <= 119090) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119091 && (row * 640 + col) <= 119626) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119627 && (row * 640 + col) <= 119627) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119628 && (row * 640 + col) <= 119635) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 119636 && (row * 640 + col) <= 119636) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119637 && (row * 640 + col) <= 119639) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 119640 && (row * 640 + col) <= 119640) color_data <= 12'b000101100000; else
        if ((row * 640 + col) >= 119641 && (row * 640 + col) <= 119642) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 119643 && (row * 640 + col) <= 119646) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119647 && (row * 640 + col) <= 119647) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 119648 && (row * 640 + col) <= 119648) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 119649 && (row * 640 + col) <= 119708) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119709 && (row * 640 + col) <= 119711) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119712 && (row * 640 + col) <= 119713) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119714 && (row * 640 + col) <= 119714) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119715 && (row * 640 + col) <= 119716) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119717 && (row * 640 + col) <= 119717) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119718 && (row * 640 + col) <= 119719) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119720 && (row * 640 + col) <= 119720) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119721 && (row * 640 + col) <= 119721) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119722 && (row * 640 + col) <= 119722) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119723 && (row * 640 + col) <= 119723) color_data <= 12'b100010110100; else
        if ((row * 640 + col) >= 119724 && (row * 640 + col) <= 119725) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 119726 && (row * 640 + col) <= 119728) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 119729 && (row * 640 + col) <= 120266) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120267 && (row * 640 + col) <= 120267) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 120268 && (row * 640 + col) <= 120269) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120270 && (row * 640 + col) <= 120270) color_data <= 12'b010010110000; else
        if ((row * 640 + col) >= 120271 && (row * 640 + col) <= 120274) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 120275 && (row * 640 + col) <= 120275) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120276 && (row * 640 + col) <= 120279) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 120280 && (row * 640 + col) <= 120280) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120281 && (row * 640 + col) <= 120284) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 120285 && (row * 640 + col) <= 120285) color_data <= 12'b011001100000; else
        if ((row * 640 + col) >= 120286 && (row * 640 + col) <= 120288) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 120289 && (row * 640 + col) <= 120289) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 120290 && (row * 640 + col) <= 120350) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120351 && (row * 640 + col) <= 120352) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120353 && (row * 640 + col) <= 120353) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 120354 && (row * 640 + col) <= 120354) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120355 && (row * 640 + col) <= 120356) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 120357 && (row * 640 + col) <= 120357) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120358 && (row * 640 + col) <= 120359) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 120360 && (row * 640 + col) <= 120361) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120362 && (row * 640 + col) <= 120364) color_data <= 12'b011010110010; else
        if ((row * 640 + col) >= 120365 && (row * 640 + col) <= 120366) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120367 && (row * 640 + col) <= 120905) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120906 && (row * 640 + col) <= 120906) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 120907 && (row * 640 + col) <= 120909) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 120910 && (row * 640 + col) <= 120915) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120916 && (row * 640 + col) <= 120918) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 120919 && (row * 640 + col) <= 120920) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 120921 && (row * 640 + col) <= 120924) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 120925 && (row * 640 + col) <= 120925) color_data <= 12'b001101100000; else
        if ((row * 640 + col) >= 120926 && (row * 640 + col) <= 120929) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 120930 && (row * 640 + col) <= 120930) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 120931 && (row * 640 + col) <= 120992) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120993 && (row * 640 + col) <= 121004) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 121005 && (row * 640 + col) <= 121545) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121546 && (row * 640 + col) <= 121546) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 121547 && (row * 640 + col) <= 121553) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 121554 && (row * 640 + col) <= 121554) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 121555 && (row * 640 + col) <= 121558) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 121559 && (row * 640 + col) <= 121559) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 121560 && (row * 640 + col) <= 121560) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 121561 && (row * 640 + col) <= 121561) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 121562 && (row * 640 + col) <= 121565) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 121566 && (row * 640 + col) <= 121566) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 121567 && (row * 640 + col) <= 121569) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 121570 && (row * 640 + col) <= 121570) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 121571 && (row * 640 + col) <= 121631) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121632 && (row * 640 + col) <= 121632) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 121633 && (row * 640 + col) <= 121635) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 121636 && (row * 640 + col) <= 121637) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 121638 && (row * 640 + col) <= 121639) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 121640 && (row * 640 + col) <= 121643) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 121644 && (row * 640 + col) <= 121645) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 121646 && (row * 640 + col) <= 122184) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122185 && (row * 640 + col) <= 122185) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 122186 && (row * 640 + col) <= 122190) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 122191 && (row * 640 + col) <= 122192) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 122193 && (row * 640 + col) <= 122193) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 122194 && (row * 640 + col) <= 122194) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 122195 && (row * 640 + col) <= 122198) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 122199 && (row * 640 + col) <= 122199) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 122200 && (row * 640 + col) <= 122200) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 122201 && (row * 640 + col) <= 122201) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 122202 && (row * 640 + col) <= 122202) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 122203 && (row * 640 + col) <= 122205) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 122206 && (row * 640 + col) <= 122206) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 122207 && (row * 640 + col) <= 122210) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 122211 && (row * 640 + col) <= 122211) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 122212 && (row * 640 + col) <= 122270) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122271 && (row * 640 + col) <= 122273) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122274 && (row * 640 + col) <= 122274) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 122275 && (row * 640 + col) <= 122276) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 122277 && (row * 640 + col) <= 122277) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 122278 && (row * 640 + col) <= 122279) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122280 && (row * 640 + col) <= 122283) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 122284 && (row * 640 + col) <= 122286) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122287 && (row * 640 + col) <= 122824) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122825 && (row * 640 + col) <= 122825) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 122826 && (row * 640 + col) <= 122826) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 122827 && (row * 640 + col) <= 122827) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 122828 && (row * 640 + col) <= 122829) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 122830 && (row * 640 + col) <= 122832) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 122833 && (row * 640 + col) <= 122833) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 122834 && (row * 640 + col) <= 122834) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 122835 && (row * 640 + col) <= 122836) color_data <= 12'b001110110000; else
        if ((row * 640 + col) >= 122837 && (row * 640 + col) <= 122838) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 122839 && (row * 640 + col) <= 122840) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 122841 && (row * 640 + col) <= 122842) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 122843 && (row * 640 + col) <= 122846) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 122847 && (row * 640 + col) <= 122850) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 122851 && (row * 640 + col) <= 122851) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 122852 && (row * 640 + col) <= 122909) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122910 && (row * 640 + col) <= 122911) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122912 && (row * 640 + col) <= 122913) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 122914 && (row * 640 + col) <= 122914) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122915 && (row * 640 + col) <= 122915) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 122916 && (row * 640 + col) <= 122916) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 122917 && (row * 640 + col) <= 122917) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122918 && (row * 640 + col) <= 122919) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 122920 && (row * 640 + col) <= 122920) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122921 && (row * 640 + col) <= 122922) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 122923 && (row * 640 + col) <= 122923) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122924 && (row * 640 + col) <= 122925) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 122926 && (row * 640 + col) <= 122927) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 122928 && (row * 640 + col) <= 123464) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123465 && (row * 640 + col) <= 123465) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 123466 && (row * 640 + col) <= 123466) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 123467 && (row * 640 + col) <= 123467) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 123468 && (row * 640 + col) <= 123468) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 123469 && (row * 640 + col) <= 123472) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 123473 && (row * 640 + col) <= 123474) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 123475 && (row * 640 + col) <= 123477) color_data <= 12'b010001100010; else
        if ((row * 640 + col) >= 123478 && (row * 640 + col) <= 123481) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 123482 && (row * 640 + col) <= 123482) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 123483 && (row * 640 + col) <= 123484) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 123485 && (row * 640 + col) <= 123490) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 123491 && (row * 640 + col) <= 123491) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 123492 && (row * 640 + col) <= 123548) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123549 && (row * 640 + col) <= 123550) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 123551 && (row * 640 + col) <= 123554) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 123555 && (row * 640 + col) <= 123556) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 123557 && (row * 640 + col) <= 123558) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 123559 && (row * 640 + col) <= 123560) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 123561 && (row * 640 + col) <= 123562) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 123563 && (row * 640 + col) <= 123566) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 123567 && (row * 640 + col) <= 123568) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 123569 && (row * 640 + col) <= 124104) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124105 && (row * 640 + col) <= 124105) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 124106 && (row * 640 + col) <= 124108) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 124109 && (row * 640 + col) <= 124111) color_data <= 12'b111111101110; else
        if ((row * 640 + col) >= 124112 && (row * 640 + col) <= 124121) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 124122 && (row * 640 + col) <= 124122) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 124123 && (row * 640 + col) <= 124125) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 124126 && (row * 640 + col) <= 124127) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 124128 && (row * 640 + col) <= 124128) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 124129 && (row * 640 + col) <= 124130) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 124131 && (row * 640 + col) <= 124131) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 124132 && (row * 640 + col) <= 124188) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124189 && (row * 640 + col) <= 124189) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124190 && (row * 640 + col) <= 124194) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 124195 && (row * 640 + col) <= 124196) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124197 && (row * 640 + col) <= 124199) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 124200 && (row * 640 + col) <= 124200) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 124201 && (row * 640 + col) <= 124202) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124203 && (row * 640 + col) <= 124207) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 124208 && (row * 640 + col) <= 124208) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124209 && (row * 640 + col) <= 124744) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124745 && (row * 640 + col) <= 124745) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 124746 && (row * 640 + col) <= 124758) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 124759 && (row * 640 + col) <= 124759) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 124760 && (row * 640 + col) <= 124761) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 124762 && (row * 640 + col) <= 124765) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 124766 && (row * 640 + col) <= 124767) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 124768 && (row * 640 + col) <= 124768) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 124769 && (row * 640 + col) <= 124770) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 124771 && (row * 640 + col) <= 124771) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 124772 && (row * 640 + col) <= 124827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124828 && (row * 640 + col) <= 124829) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124830 && (row * 640 + col) <= 124833) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 124834 && (row * 640 + col) <= 124834) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124835 && (row * 640 + col) <= 124835) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 124836 && (row * 640 + col) <= 124836) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 124837 && (row * 640 + col) <= 124837) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124838 && (row * 640 + col) <= 124839) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 124840 && (row * 640 + col) <= 124840) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124841 && (row * 640 + col) <= 124842) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 124843 && (row * 640 + col) <= 124843) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124844 && (row * 640 + col) <= 124847) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 124848 && (row * 640 + col) <= 124849) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 124850 && (row * 640 + col) <= 125384) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125385 && (row * 640 + col) <= 125385) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 125386 && (row * 640 + col) <= 125390) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 125391 && (row * 640 + col) <= 125391) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 125392 && (row * 640 + col) <= 125398) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 125399 && (row * 640 + col) <= 125399) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 125400 && (row * 640 + col) <= 125401) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 125402 && (row * 640 + col) <= 125406) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 125407 && (row * 640 + col) <= 125410) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 125411 && (row * 640 + col) <= 125411) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 125412 && (row * 640 + col) <= 125467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125468 && (row * 640 + col) <= 125468) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 125469 && (row * 640 + col) <= 125469) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 125470 && (row * 640 + col) <= 125470) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 125471 && (row * 640 + col) <= 125472) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 125473 && (row * 640 + col) <= 125473) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 125474 && (row * 640 + col) <= 125474) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 125475 && (row * 640 + col) <= 125477) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 125478 && (row * 640 + col) <= 125479) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 125480 && (row * 640 + col) <= 125480) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 125481 && (row * 640 + col) <= 125483) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 125484 && (row * 640 + col) <= 125484) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 125485 && (row * 640 + col) <= 125486) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 125487 && (row * 640 + col) <= 125487) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 125488 && (row * 640 + col) <= 125488) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 125489 && (row * 640 + col) <= 125489) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 125490 && (row * 640 + col) <= 126024) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126025 && (row * 640 + col) <= 126025) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 126026 && (row * 640 + col) <= 126030) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 126031 && (row * 640 + col) <= 126031) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 126032 && (row * 640 + col) <= 126041) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 126042 && (row * 640 + col) <= 126046) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 126047 && (row * 640 + col) <= 126050) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 126051 && (row * 640 + col) <= 126051) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 126052 && (row * 640 + col) <= 126107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126108 && (row * 640 + col) <= 126108) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126109 && (row * 640 + col) <= 126109) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 126110 && (row * 640 + col) <= 126110) color_data <= 12'b111111111100; else
        if ((row * 640 + col) >= 126111 && (row * 640 + col) <= 126112) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126113 && (row * 640 + col) <= 126117) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 126118 && (row * 640 + col) <= 126119) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126120 && (row * 640 + col) <= 126121) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 126122 && (row * 640 + col) <= 126124) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 126125 && (row * 640 + col) <= 126126) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126127 && (row * 640 + col) <= 126128) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 126129 && (row * 640 + col) <= 126129) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126130 && (row * 640 + col) <= 126664) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126665 && (row * 640 + col) <= 126665) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 126666 && (row * 640 + col) <= 126666) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 126667 && (row * 640 + col) <= 126667) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 126668 && (row * 640 + col) <= 126675) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 126676 && (row * 640 + col) <= 126676) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 126677 && (row * 640 + col) <= 126680) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 126681 && (row * 640 + col) <= 126682) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 126683 && (row * 640 + col) <= 126683) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 126684 && (row * 640 + col) <= 126686) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 126687 && (row * 640 + col) <= 126689) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 126690 && (row * 640 + col) <= 126690) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 126691 && (row * 640 + col) <= 126691) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 126692 && (row * 640 + col) <= 126747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126748 && (row * 640 + col) <= 126748) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126749 && (row * 640 + col) <= 126750) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 126751 && (row * 640 + col) <= 126752) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126753 && (row * 640 + col) <= 126755) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 126756 && (row * 640 + col) <= 126757) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126758 && (row * 640 + col) <= 126759) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 126760 && (row * 640 + col) <= 126761) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126762 && (row * 640 + col) <= 126764) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 126765 && (row * 640 + col) <= 126766) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126767 && (row * 640 + col) <= 126768) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 126769 && (row * 640 + col) <= 126769) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 126770 && (row * 640 + col) <= 127304) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127305 && (row * 640 + col) <= 127305) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 127306 && (row * 640 + col) <= 127306) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 127307 && (row * 640 + col) <= 127307) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 127308 && (row * 640 + col) <= 127315) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 127316 && (row * 640 + col) <= 127316) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 127317 && (row * 640 + col) <= 127320) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 127321 && (row * 640 + col) <= 127322) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 127323 && (row * 640 + col) <= 127323) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 127324 && (row * 640 + col) <= 127326) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 127327 && (row * 640 + col) <= 127329) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 127330 && (row * 640 + col) <= 127330) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 127331 && (row * 640 + col) <= 127331) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 127332 && (row * 640 + col) <= 127387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127388 && (row * 640 + col) <= 127388) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127389 && (row * 640 + col) <= 127389) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 127390 && (row * 640 + col) <= 127390) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127391 && (row * 640 + col) <= 127392) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 127393 && (row * 640 + col) <= 127393) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127394 && (row * 640 + col) <= 127394) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 127395 && (row * 640 + col) <= 127395) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127396 && (row * 640 + col) <= 127401) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 127402 && (row * 640 + col) <= 127402) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127403 && (row * 640 + col) <= 127403) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 127404 && (row * 640 + col) <= 127404) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127405 && (row * 640 + col) <= 127406) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 127407 && (row * 640 + col) <= 127407) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127408 && (row * 640 + col) <= 127408) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 127409 && (row * 640 + col) <= 127409) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 127410 && (row * 640 + col) <= 127944) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127945 && (row * 640 + col) <= 127945) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 127946 && (row * 640 + col) <= 127958) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 127959 && (row * 640 + col) <= 127965) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 127966 && (row * 640 + col) <= 127970) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 127971 && (row * 640 + col) <= 127971) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 127972 && (row * 640 + col) <= 128027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128028 && (row * 640 + col) <= 128029) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128030 && (row * 640 + col) <= 128033) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 128034 && (row * 640 + col) <= 128034) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128035 && (row * 640 + col) <= 128040) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 128041 && (row * 640 + col) <= 128042) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 128043 && (row * 640 + col) <= 128043) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128044 && (row * 640 + col) <= 128047) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 128048 && (row * 640 + col) <= 128049) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128050 && (row * 640 + col) <= 128585) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128586 && (row * 640 + col) <= 128586) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 128587 && (row * 640 + col) <= 128597) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 128598 && (row * 640 + col) <= 128605) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 128606 && (row * 640 + col) <= 128609) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 128610 && (row * 640 + col) <= 128610) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 128611 && (row * 640 + col) <= 128667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128668 && (row * 640 + col) <= 128668) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128669 && (row * 640 + col) <= 128673) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 128674 && (row * 640 + col) <= 128674) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128675 && (row * 640 + col) <= 128680) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 128681 && (row * 640 + col) <= 128682) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 128683 && (row * 640 + col) <= 128683) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128684 && (row * 640 + col) <= 128688) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 128689 && (row * 640 + col) <= 128689) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 128690 && (row * 640 + col) <= 129226) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129227 && (row * 640 + col) <= 129227) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 129228 && (row * 640 + col) <= 129229) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 129230 && (row * 640 + col) <= 129230) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129231 && (row * 640 + col) <= 129233) color_data <= 12'b111100100000; else
        if ((row * 640 + col) >= 129234 && (row * 640 + col) <= 129238) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 129239 && (row * 640 + col) <= 129239) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129240 && (row * 640 + col) <= 129244) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 129245 && (row * 640 + col) <= 129246) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 129247 && (row * 640 + col) <= 129247) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129248 && (row * 640 + col) <= 129248) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 129249 && (row * 640 + col) <= 129249) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 129250 && (row * 640 + col) <= 129307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129308 && (row * 640 + col) <= 129308) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129309 && (row * 640 + col) <= 129312) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 129313 && (row * 640 + col) <= 129313) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129314 && (row * 640 + col) <= 129314) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 129315 && (row * 640 + col) <= 129315) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129316 && (row * 640 + col) <= 129319) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 129320 && (row * 640 + col) <= 129321) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 129322 && (row * 640 + col) <= 129322) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129323 && (row * 640 + col) <= 129323) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 129324 && (row * 640 + col) <= 129324) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129325 && (row * 640 + col) <= 129328) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 129329 && (row * 640 + col) <= 129329) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129330 && (row * 640 + col) <= 129866) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129867 && (row * 640 + col) <= 129867) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 129868 && (row * 640 + col) <= 129868) color_data <= 12'b101000010001; else
        if ((row * 640 + col) >= 129869 && (row * 640 + col) <= 129869) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 129870 && (row * 640 + col) <= 129870) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129871 && (row * 640 + col) <= 129874) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 129875 && (row * 640 + col) <= 129875) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129876 && (row * 640 + col) <= 129878) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 129879 && (row * 640 + col) <= 129879) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129880 && (row * 640 + col) <= 129882) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 129883 && (row * 640 + col) <= 129883) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129884 && (row * 640 + col) <= 129886) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 129887 && (row * 640 + col) <= 129887) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 129888 && (row * 640 + col) <= 129888) color_data <= 12'b100100000000; else
        if ((row * 640 + col) >= 129889 && (row * 640 + col) <= 129889) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 129890 && (row * 640 + col) <= 129947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129948 && (row * 640 + col) <= 129949) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129950 && (row * 640 + col) <= 129951) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 129952 && (row * 640 + col) <= 129952) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129953 && (row * 640 + col) <= 129955) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 129956 && (row * 640 + col) <= 129957) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129958 && (row * 640 + col) <= 129958) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 129959 && (row * 640 + col) <= 129959) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 129960 && (row * 640 + col) <= 129961) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129962 && (row * 640 + col) <= 129964) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 129965 && (row * 640 + col) <= 129965) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129966 && (row * 640 + col) <= 129967) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 129968 && (row * 640 + col) <= 129969) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 129970 && (row * 640 + col) <= 130507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130508 && (row * 640 + col) <= 130508) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 130509 && (row * 640 + col) <= 130514) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 130515 && (row * 640 + col) <= 130515) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 130516 && (row * 640 + col) <= 130522) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 130523 && (row * 640 + col) <= 130523) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 130524 && (row * 640 + col) <= 130527) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 130528 && (row * 640 + col) <= 130528) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 130529 && (row * 640 + col) <= 130587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130588 && (row * 640 + col) <= 130588) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 130589 && (row * 640 + col) <= 130589) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 130590 && (row * 640 + col) <= 130591) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 130592 && (row * 640 + col) <= 130597) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 130598 && (row * 640 + col) <= 130599) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 130600 && (row * 640 + col) <= 130605) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 130606 && (row * 640 + col) <= 130607) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 130608 && (row * 640 + col) <= 130608) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 130609 && (row * 640 + col) <= 130609) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 130610 && (row * 640 + col) <= 131148) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131149 && (row * 640 + col) <= 131149) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 131150 && (row * 640 + col) <= 131161) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 131162 && (row * 640 + col) <= 131166) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 131167 && (row * 640 + col) <= 131167) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 131168 && (row * 640 + col) <= 131227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131228 && (row * 640 + col) <= 131228) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131229 && (row * 640 + col) <= 131229) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 131230 && (row * 640 + col) <= 131231) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131232 && (row * 640 + col) <= 131237) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 131238 && (row * 640 + col) <= 131239) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131240 && (row * 640 + col) <= 131245) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 131246 && (row * 640 + col) <= 131247) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131248 && (row * 640 + col) <= 131248) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 131249 && (row * 640 + col) <= 131249) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131250 && (row * 640 + col) <= 131789) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131790 && (row * 640 + col) <= 131790) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 131791 && (row * 640 + col) <= 131791) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 131792 && (row * 640 + col) <= 131800) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 131801 && (row * 640 + col) <= 131805) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 131806 && (row * 640 + col) <= 131806) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 131807 && (row * 640 + col) <= 131867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131868 && (row * 640 + col) <= 131869) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131870 && (row * 640 + col) <= 131871) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 131872 && (row * 640 + col) <= 131872) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131873 && (row * 640 + col) <= 131876) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 131877 && (row * 640 + col) <= 131877) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 131878 && (row * 640 + col) <= 131879) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131880 && (row * 640 + col) <= 131884) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 131885 && (row * 640 + col) <= 131885) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131886 && (row * 640 + col) <= 131887) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 131888 && (row * 640 + col) <= 131889) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 131890 && (row * 640 + col) <= 132430) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132431 && (row * 640 + col) <= 132431) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 132432 && (row * 640 + col) <= 132432) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 132433 && (row * 640 + col) <= 132436) color_data <= 12'b111000010000; else
        if ((row * 640 + col) >= 132437 && (row * 640 + col) <= 132441) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 132442 && (row * 640 + col) <= 132442) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 132443 && (row * 640 + col) <= 132444) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 132445 && (row * 640 + col) <= 132445) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 132446 && (row * 640 + col) <= 132507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132508 && (row * 640 + col) <= 132508) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 132509 && (row * 640 + col) <= 132510) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 132511 && (row * 640 + col) <= 132512) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 132513 && (row * 640 + col) <= 132513) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 132514 && (row * 640 + col) <= 132515) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 132516 && (row * 640 + col) <= 132517) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 132518 && (row * 640 + col) <= 132519) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 132520 && (row * 640 + col) <= 132521) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 132522 && (row * 640 + col) <= 132523) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 132524 && (row * 640 + col) <= 132524) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 132525 && (row * 640 + col) <= 132528) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 132529 && (row * 640 + col) <= 132529) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 132530 && (row * 640 + col) <= 133071) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133072 && (row * 640 + col) <= 133072) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 133073 && (row * 640 + col) <= 133073) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 133074 && (row * 640 + col) <= 133081) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 133082 && (row * 640 + col) <= 133082) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 133083 && (row * 640 + col) <= 133083) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 133084 && (row * 640 + col) <= 133084) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 133085 && (row * 640 + col) <= 133147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133148 && (row * 640 + col) <= 133149) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133150 && (row * 640 + col) <= 133151) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 133152 && (row * 640 + col) <= 133153) color_data <= 12'b111111110011; else
        if ((row * 640 + col) >= 133154 && (row * 640 + col) <= 133155) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133156 && (row * 640 + col) <= 133161) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 133162 && (row * 640 + col) <= 133163) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133164 && (row * 640 + col) <= 133167) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 133168 && (row * 640 + col) <= 133169) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133170 && (row * 640 + col) <= 133712) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133713 && (row * 640 + col) <= 133713) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 133714 && (row * 640 + col) <= 133716) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 133717 && (row * 640 + col) <= 133717) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 133718 && (row * 640 + col) <= 133722) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 133723 && (row * 640 + col) <= 133723) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 133724 && (row * 640 + col) <= 133788) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133789 && (row * 640 + col) <= 133789) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133790 && (row * 640 + col) <= 133793) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 133794 && (row * 640 + col) <= 133795) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133796 && (row * 640 + col) <= 133801) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 133802 && (row * 640 + col) <= 133803) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133804 && (row * 640 + col) <= 133807) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 133808 && (row * 640 + col) <= 133808) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 133809 && (row * 640 + col) <= 134353) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134354 && (row * 640 + col) <= 134354) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 134355 && (row * 640 + col) <= 134356) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 134357 && (row * 640 + col) <= 134357) color_data <= 12'b111110110000; else
        if ((row * 640 + col) >= 134358 && (row * 640 + col) <= 134361) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 134362 && (row * 640 + col) <= 134362) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 134363 && (row * 640 + col) <= 134428) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134429 && (row * 640 + col) <= 134430) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 134431 && (row * 640 + col) <= 134432) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 134433 && (row * 640 + col) <= 134433) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 134434 && (row * 640 + col) <= 134435) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 134436 && (row * 640 + col) <= 134436) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 134437 && (row * 640 + col) <= 134440) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 134441 && (row * 640 + col) <= 134441) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 134442 && (row * 640 + col) <= 134443) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 134444 && (row * 640 + col) <= 134444) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 134445 && (row * 640 + col) <= 134446) color_data <= 12'b111011000000; else
        if ((row * 640 + col) >= 134447 && (row * 640 + col) <= 134448) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 134449 && (row * 640 + col) <= 134994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134995 && (row * 640 + col) <= 134996) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 134997 && (row * 640 + col) <= 134999) color_data <= 12'b110000000000; else
        if ((row * 640 + col) >= 135000 && (row * 640 + col) <= 135001) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 135002 && (row * 640 + col) <= 135069) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135070 && (row * 640 + col) <= 135087) color_data <= 12'b100101100000; else
        if ((row * 640 + col) >= 135088 && (row * 640 + col) <= 135636) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135637 && (row * 640 + col) <= 135639) color_data <= 12'b100100010000; else
        if ((row * 640 + col) >= 135640 && (row * 640 + col) <= 145038) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145039 && (row * 640 + col) <= 145041) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 145042 && (row * 640 + col) <= 145678) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145679 && (row * 640 + col) <= 145681) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 145682 && (row * 640 + col) <= 146318) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 146319 && (row * 640 + col) <= 146321) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 146322 && (row * 640 + col) <= 146958) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 146959 && (row * 640 + col) <= 146961) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 146962 && (row * 640 + col) <= 147598) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 147599 && (row * 640 + col) <= 147601) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 147602 && (row * 640 + col) <= 148238) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 148239 && (row * 640 + col) <= 148241) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 148242 && (row * 640 + col) <= 148479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 148480 && (row * 640 + col) <= 148485) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 148486 && (row * 640 + col) <= 148878) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 148879 && (row * 640 + col) <= 148881) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 148882 && (row * 640 + col) <= 149119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149120 && (row * 640 + col) <= 149125) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 149126 && (row * 640 + col) <= 149518) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149519 && (row * 640 + col) <= 149521) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149522 && (row * 640 + col) <= 149759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149760 && (row * 640 + col) <= 149766) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 149767 && (row * 640 + col) <= 149970) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149971 && (row * 640 + col) <= 149980) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 149981 && (row * 640 + col) <= 150158) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 150159 && (row * 640 + col) <= 150161) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150162 && (row * 640 + col) <= 150399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 150400 && (row * 640 + col) <= 150419) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 150420 && (row * 640 + col) <= 150607) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 150608 && (row * 640 + col) <= 150623) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 150624 && (row * 640 + col) <= 150798) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 150799 && (row * 640 + col) <= 150801) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150802 && (row * 640 + col) <= 151039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151040 && (row * 640 + col) <= 151059) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151060 && (row * 640 + col) <= 151245) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151246 && (row * 640 + col) <= 151251) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 151252 && (row * 640 + col) <= 151259) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 151260 && (row * 640 + col) <= 151265) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 151266 && (row * 640 + col) <= 151438) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151439 && (row * 640 + col) <= 151441) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151442 && (row * 640 + col) <= 151679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151680 && (row * 640 + col) <= 151704) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151705 && (row * 640 + col) <= 151884) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151885 && (row * 640 + col) <= 151888) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 151889 && (row * 640 + col) <= 151902) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 151903 && (row * 640 + col) <= 151906) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 151907 && (row * 640 + col) <= 152078) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152079 && (row * 640 + col) <= 152081) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152082 && (row * 640 + col) <= 152319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152320 && (row * 640 + col) <= 152345) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 152346 && (row * 640 + col) <= 152523) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152524 && (row * 640 + col) <= 152526) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 152527 && (row * 640 + col) <= 152544) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 152545 && (row * 640 + col) <= 152547) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 152548 && (row * 640 + col) <= 152718) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152719 && (row * 640 + col) <= 152721) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152722 && (row * 640 + col) <= 152959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152960 && (row * 640 + col) <= 152985) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 152986 && (row * 640 + col) <= 153162) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153163 && (row * 640 + col) <= 153165) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 153166 && (row * 640 + col) <= 153185) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 153186 && (row * 640 + col) <= 153188) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 153189 && (row * 640 + col) <= 153358) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153359 && (row * 640 + col) <= 153361) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153362 && (row * 640 + col) <= 153599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153600 && (row * 640 + col) <= 153627) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 153628 && (row * 640 + col) <= 153801) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153802 && (row * 640 + col) <= 153804) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 153805 && (row * 640 + col) <= 153826) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 153827 && (row * 640 + col) <= 153829) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 153830 && (row * 640 + col) <= 153998) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153999 && (row * 640 + col) <= 154001) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154002 && (row * 640 + col) <= 154239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154240 && (row * 640 + col) <= 154270) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 154271 && (row * 640 + col) <= 154440) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154441 && (row * 640 + col) <= 154443) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 154444 && (row * 640 + col) <= 154467) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 154468 && (row * 640 + col) <= 154470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 154471 && (row * 640 + col) <= 154638) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154639 && (row * 640 + col) <= 154641) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154642 && (row * 640 + col) <= 154879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154880 && (row * 640 + col) <= 154911) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 154912 && (row * 640 + col) <= 155079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155080 && (row * 640 + col) <= 155082) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155083 && (row * 640 + col) <= 155108) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 155109 && (row * 640 + col) <= 155111) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155112 && (row * 640 + col) <= 155278) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155279 && (row * 640 + col) <= 155281) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155282 && (row * 640 + col) <= 155519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155520 && (row * 640 + col) <= 155552) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155553 && (row * 640 + col) <= 155718) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155719 && (row * 640 + col) <= 155721) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155722 && (row * 640 + col) <= 155749) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 155750 && (row * 640 + col) <= 155752) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155753 && (row * 640 + col) <= 155794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155795 && (row * 640 + col) <= 155809) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155810 && (row * 640 + col) <= 155812) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155813 && (row * 640 + col) <= 155824) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155825 && (row * 640 + col) <= 155827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155828 && (row * 640 + col) <= 155842) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155843 && (row * 640 + col) <= 155845) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155846 && (row * 640 + col) <= 155860) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155861 && (row * 640 + col) <= 155863) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155864 && (row * 640 + col) <= 155875) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155876 && (row * 640 + col) <= 155884) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155885 && (row * 640 + col) <= 155899) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155900 && (row * 640 + col) <= 155902) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155903 && (row * 640 + col) <= 155917) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155918 && (row * 640 + col) <= 155918) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155919 && (row * 640 + col) <= 155920) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155921 && (row * 640 + col) <= 155926) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155927 && (row * 640 + col) <= 155935) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155936 && (row * 640 + col) <= 155941) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155942 && (row * 640 + col) <= 155944) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155945 && (row * 640 + col) <= 155959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155960 && (row * 640 + col) <= 155962) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155963 && (row * 640 + col) <= 155968) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 155969 && (row * 640 + col) <= 156159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156160 && (row * 640 + col) <= 156193) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 156194 && (row * 640 + col) <= 156358) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156359 && (row * 640 + col) <= 156360) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156361 && (row * 640 + col) <= 156390) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 156391 && (row * 640 + col) <= 156392) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156393 && (row * 640 + col) <= 156434) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156435 && (row * 640 + col) <= 156449) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156450 && (row * 640 + col) <= 156452) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156453 && (row * 640 + col) <= 156464) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156465 && (row * 640 + col) <= 156467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156468 && (row * 640 + col) <= 156482) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156483 && (row * 640 + col) <= 156485) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156486 && (row * 640 + col) <= 156500) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156501 && (row * 640 + col) <= 156503) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156504 && (row * 640 + col) <= 156515) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156516 && (row * 640 + col) <= 156524) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156525 && (row * 640 + col) <= 156539) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156540 && (row * 640 + col) <= 156542) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156543 && (row * 640 + col) <= 156557) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156558 && (row * 640 + col) <= 156558) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156559 && (row * 640 + col) <= 156560) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156561 && (row * 640 + col) <= 156566) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156567 && (row * 640 + col) <= 156575) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156576 && (row * 640 + col) <= 156581) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156582 && (row * 640 + col) <= 156584) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156585 && (row * 640 + col) <= 156599) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156600 && (row * 640 + col) <= 156602) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156603 && (row * 640 + col) <= 156608) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 156609 && (row * 640 + col) <= 156799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156800 && (row * 640 + col) <= 156834) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 156835 && (row * 640 + col) <= 156997) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156998 && (row * 640 + col) <= 157000) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157001 && (row * 640 + col) <= 157030) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 157031 && (row * 640 + col) <= 157033) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157034 && (row * 640 + col) <= 157074) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157075 && (row * 640 + col) <= 157089) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157090 && (row * 640 + col) <= 157092) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157093 && (row * 640 + col) <= 157104) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157105 && (row * 640 + col) <= 157107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157108 && (row * 640 + col) <= 157122) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157123 && (row * 640 + col) <= 157125) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157126 && (row * 640 + col) <= 157140) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157141 && (row * 640 + col) <= 157143) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157144 && (row * 640 + col) <= 157155) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157156 && (row * 640 + col) <= 157164) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157165 && (row * 640 + col) <= 157179) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157180 && (row * 640 + col) <= 157182) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157183 && (row * 640 + col) <= 157197) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157198 && (row * 640 + col) <= 157198) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157199 && (row * 640 + col) <= 157200) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157201 && (row * 640 + col) <= 157206) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157207 && (row * 640 + col) <= 157215) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157216 && (row * 640 + col) <= 157221) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157222 && (row * 640 + col) <= 157224) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157225 && (row * 640 + col) <= 157239) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157240 && (row * 640 + col) <= 157242) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157243 && (row * 640 + col) <= 157248) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157249 && (row * 640 + col) <= 157439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157440 && (row * 640 + col) <= 157493) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157494 && (row * 640 + col) <= 157637) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157638 && (row * 640 + col) <= 157639) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157640 && (row * 640 + col) <= 157671) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 157672 && (row * 640 + col) <= 157673) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157674 && (row * 640 + col) <= 157691) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157692 && (row * 640 + col) <= 157695) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157696 && (row * 640 + col) <= 157714) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157715 && (row * 640 + col) <= 157720) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157721 && (row * 640 + col) <= 157723) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157724 && (row * 640 + col) <= 157729) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157730 && (row * 640 + col) <= 157735) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157736 && (row * 640 + col) <= 157741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157742 && (row * 640 + col) <= 157747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157748 && (row * 640 + col) <= 157753) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157754 && (row * 640 + col) <= 157756) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157757 && (row * 640 + col) <= 157762) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157763 && (row * 640 + col) <= 157765) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157766 && (row * 640 + col) <= 157771) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157772 && (row * 640 + col) <= 157774) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157775 && (row * 640 + col) <= 157780) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157781 && (row * 640 + col) <= 157786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157787 && (row * 640 + col) <= 157792) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157793 && (row * 640 + col) <= 157804) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157805 && (row * 640 + col) <= 157810) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157811 && (row * 640 + col) <= 157813) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157814 && (row * 640 + col) <= 157819) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157820 && (row * 640 + col) <= 157822) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157823 && (row * 640 + col) <= 157828) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157829 && (row * 640 + col) <= 157831) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157832 && (row * 640 + col) <= 157837) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157838 && (row * 640 + col) <= 157838) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157839 && (row * 640 + col) <= 157840) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157841 && (row * 640 + col) <= 157849) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157850 && (row * 640 + col) <= 157852) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157853 && (row * 640 + col) <= 157861) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157862 && (row * 640 + col) <= 157864) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157865 && (row * 640 + col) <= 157870) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157871 && (row * 640 + col) <= 157873) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157874 && (row * 640 + col) <= 157879) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157880 && (row * 640 + col) <= 157882) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157883 && (row * 640 + col) <= 157888) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 157889 && (row * 640 + col) <= 158079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158080 && (row * 640 + col) <= 158133) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 158134 && (row * 640 + col) <= 158277) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158278 && (row * 640 + col) <= 158279) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158280 && (row * 640 + col) <= 158311) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 158312 && (row * 640 + col) <= 158313) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158314 && (row * 640 + col) <= 158331) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158332 && (row * 640 + col) <= 158335) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158336 && (row * 640 + col) <= 158354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158355 && (row * 640 + col) <= 158360) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158361 && (row * 640 + col) <= 158363) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158364 && (row * 640 + col) <= 158369) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158370 && (row * 640 + col) <= 158375) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158376 && (row * 640 + col) <= 158381) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158382 && (row * 640 + col) <= 158387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158388 && (row * 640 + col) <= 158393) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158394 && (row * 640 + col) <= 158396) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158397 && (row * 640 + col) <= 158402) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158403 && (row * 640 + col) <= 158405) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158406 && (row * 640 + col) <= 158411) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158412 && (row * 640 + col) <= 158414) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158415 && (row * 640 + col) <= 158420) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158421 && (row * 640 + col) <= 158426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158427 && (row * 640 + col) <= 158432) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158433 && (row * 640 + col) <= 158444) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158445 && (row * 640 + col) <= 158450) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158451 && (row * 640 + col) <= 158453) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158454 && (row * 640 + col) <= 158459) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158460 && (row * 640 + col) <= 158462) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158463 && (row * 640 + col) <= 158468) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158469 && (row * 640 + col) <= 158471) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158472 && (row * 640 + col) <= 158477) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158478 && (row * 640 + col) <= 158478) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158479 && (row * 640 + col) <= 158480) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158481 && (row * 640 + col) <= 158489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158490 && (row * 640 + col) <= 158492) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158493 && (row * 640 + col) <= 158501) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158502 && (row * 640 + col) <= 158504) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158505 && (row * 640 + col) <= 158510) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158511 && (row * 640 + col) <= 158513) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158514 && (row * 640 + col) <= 158519) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158520 && (row * 640 + col) <= 158522) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158523 && (row * 640 + col) <= 158528) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158529 && (row * 640 + col) <= 158719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158720 && (row * 640 + col) <= 158774) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 158775 && (row * 640 + col) <= 158916) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158917 && (row * 640 + col) <= 158919) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158920 && (row * 640 + col) <= 158951) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 158952 && (row * 640 + col) <= 158954) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158955 && (row * 640 + col) <= 158971) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158972 && (row * 640 + col) <= 158975) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 158976 && (row * 640 + col) <= 158994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158995 && (row * 640 + col) <= 159000) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159001 && (row * 640 + col) <= 159003) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159004 && (row * 640 + col) <= 159009) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159010 && (row * 640 + col) <= 159015) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159016 && (row * 640 + col) <= 159021) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159022 && (row * 640 + col) <= 159027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159028 && (row * 640 + col) <= 159033) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159034 && (row * 640 + col) <= 159036) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159037 && (row * 640 + col) <= 159042) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159043 && (row * 640 + col) <= 159045) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159046 && (row * 640 + col) <= 159051) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159052 && (row * 640 + col) <= 159054) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159055 && (row * 640 + col) <= 159060) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159061 && (row * 640 + col) <= 159066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159067 && (row * 640 + col) <= 159072) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159073 && (row * 640 + col) <= 159084) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159085 && (row * 640 + col) <= 159090) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159091 && (row * 640 + col) <= 159093) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159094 && (row * 640 + col) <= 159099) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159100 && (row * 640 + col) <= 159102) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159103 && (row * 640 + col) <= 159108) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159109 && (row * 640 + col) <= 159111) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159112 && (row * 640 + col) <= 159117) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159118 && (row * 640 + col) <= 159118) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159119 && (row * 640 + col) <= 159120) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159121 && (row * 640 + col) <= 159129) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159130 && (row * 640 + col) <= 159132) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159133 && (row * 640 + col) <= 159141) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159142 && (row * 640 + col) <= 159144) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159145 && (row * 640 + col) <= 159150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159151 && (row * 640 + col) <= 159153) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159154 && (row * 640 + col) <= 159159) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159160 && (row * 640 + col) <= 159162) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159163 && (row * 640 + col) <= 159168) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159169 && (row * 640 + col) <= 159359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159360 && (row * 640 + col) <= 159419) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 159420 && (row * 640 + col) <= 159556) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159557 && (row * 640 + col) <= 159558) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159559 && (row * 640 + col) <= 159562) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 159563 && (row * 640 + col) <= 159567) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 159568 && (row * 640 + col) <= 159568) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 159569 && (row * 640 + col) <= 159572) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 159573 && (row * 640 + col) <= 159573) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 159574 && (row * 640 + col) <= 159578) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 159579 && (row * 640 + col) <= 159579) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 159580 && (row * 640 + col) <= 159584) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 159585 && (row * 640 + col) <= 159585) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 159586 && (row * 640 + col) <= 159589) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 159590 && (row * 640 + col) <= 159592) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 159593 && (row * 640 + col) <= 159594) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159595 && (row * 640 + col) <= 159611) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159612 && (row * 640 + col) <= 159615) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159616 && (row * 640 + col) <= 159634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159635 && (row * 640 + col) <= 159640) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159641 && (row * 640 + col) <= 159655) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159656 && (row * 640 + col) <= 159661) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159662 && (row * 640 + col) <= 159667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159668 && (row * 640 + col) <= 159673) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159674 && (row * 640 + col) <= 159676) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159677 && (row * 640 + col) <= 159682) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159683 && (row * 640 + col) <= 159685) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159686 && (row * 640 + col) <= 159691) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159692 && (row * 640 + col) <= 159694) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159695 && (row * 640 + col) <= 159700) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159701 && (row * 640 + col) <= 159706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159707 && (row * 640 + col) <= 159712) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159713 && (row * 640 + col) <= 159724) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159725 && (row * 640 + col) <= 159730) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159731 && (row * 640 + col) <= 159742) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159743 && (row * 640 + col) <= 159748) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159749 && (row * 640 + col) <= 159751) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159752 && (row * 640 + col) <= 159757) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159758 && (row * 640 + col) <= 159758) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159759 && (row * 640 + col) <= 159760) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159761 && (row * 640 + col) <= 159781) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159782 && (row * 640 + col) <= 159784) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159785 && (row * 640 + col) <= 159790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159791 && (row * 640 + col) <= 159802) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159803 && (row * 640 + col) <= 159808) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 159809 && (row * 640 + col) <= 159999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160000 && (row * 640 + col) <= 160059) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160060 && (row * 640 + col) <= 160196) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160197 && (row * 640 + col) <= 160198) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160199 && (row * 640 + col) <= 160202) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160203 && (row * 640 + col) <= 160204) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160205 && (row * 640 + col) <= 160205) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160206 && (row * 640 + col) <= 160207) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160208 && (row * 640 + col) <= 160209) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160210 && (row * 640 + col) <= 160211) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160212 && (row * 640 + col) <= 160213) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160214 && (row * 640 + col) <= 160215) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160216 && (row * 640 + col) <= 160216) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160217 && (row * 640 + col) <= 160218) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160219 && (row * 640 + col) <= 160219) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160220 && (row * 640 + col) <= 160221) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160222 && (row * 640 + col) <= 160222) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160223 && (row * 640 + col) <= 160224) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160225 && (row * 640 + col) <= 160226) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160227 && (row * 640 + col) <= 160228) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160229 && (row * 640 + col) <= 160232) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160233 && (row * 640 + col) <= 160234) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160235 && (row * 640 + col) <= 160274) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160275 && (row * 640 + col) <= 160280) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160281 && (row * 640 + col) <= 160295) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160296 && (row * 640 + col) <= 160301) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160302 && (row * 640 + col) <= 160307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160308 && (row * 640 + col) <= 160313) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160314 && (row * 640 + col) <= 160316) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160317 && (row * 640 + col) <= 160322) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160323 && (row * 640 + col) <= 160325) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160326 && (row * 640 + col) <= 160331) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160332 && (row * 640 + col) <= 160334) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160335 && (row * 640 + col) <= 160340) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160341 && (row * 640 + col) <= 160346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160347 && (row * 640 + col) <= 160352) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160353 && (row * 640 + col) <= 160364) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160365 && (row * 640 + col) <= 160370) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160371 && (row * 640 + col) <= 160382) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160383 && (row * 640 + col) <= 160388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160389 && (row * 640 + col) <= 160391) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160392 && (row * 640 + col) <= 160397) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160398 && (row * 640 + col) <= 160398) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160399 && (row * 640 + col) <= 160400) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160401 && (row * 640 + col) <= 160421) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160422 && (row * 640 + col) <= 160424) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160425 && (row * 640 + col) <= 160430) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160431 && (row * 640 + col) <= 160442) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160443 && (row * 640 + col) <= 160448) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160449 && (row * 640 + col) <= 160639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160640 && (row * 640 + col) <= 160699) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160700 && (row * 640 + col) <= 160836) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160837 && (row * 640 + col) <= 160838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160839 && (row * 640 + col) <= 160842) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160843 && (row * 640 + col) <= 160844) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160845 && (row * 640 + col) <= 160849) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160850 && (row * 640 + col) <= 160851) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160852 && (row * 640 + col) <= 160853) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160854 && (row * 640 + col) <= 160855) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160856 && (row * 640 + col) <= 160856) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160857 && (row * 640 + col) <= 160858) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160859 && (row * 640 + col) <= 160859) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160860 && (row * 640 + col) <= 160861) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160862 && (row * 640 + col) <= 160862) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160863 && (row * 640 + col) <= 160864) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160865 && (row * 640 + col) <= 160866) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160867 && (row * 640 + col) <= 160868) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 160869 && (row * 640 + col) <= 160872) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 160873 && (row * 640 + col) <= 160874) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160875 && (row * 640 + col) <= 160914) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160915 && (row * 640 + col) <= 160920) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160921 && (row * 640 + col) <= 160935) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160936 && (row * 640 + col) <= 160941) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160942 && (row * 640 + col) <= 160947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160948 && (row * 640 + col) <= 160953) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160954 && (row * 640 + col) <= 160956) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160957 && (row * 640 + col) <= 160962) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160963 && (row * 640 + col) <= 160965) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160966 && (row * 640 + col) <= 160971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160972 && (row * 640 + col) <= 160974) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160975 && (row * 640 + col) <= 160980) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160981 && (row * 640 + col) <= 160986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160987 && (row * 640 + col) <= 160992) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 160993 && (row * 640 + col) <= 161004) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161005 && (row * 640 + col) <= 161010) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161011 && (row * 640 + col) <= 161022) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161023 && (row * 640 + col) <= 161028) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161029 && (row * 640 + col) <= 161031) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161032 && (row * 640 + col) <= 161037) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161038 && (row * 640 + col) <= 161038) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161039 && (row * 640 + col) <= 161040) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161041 && (row * 640 + col) <= 161061) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161062 && (row * 640 + col) <= 161064) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161065 && (row * 640 + col) <= 161070) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161071 && (row * 640 + col) <= 161082) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161083 && (row * 640 + col) <= 161088) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161089 && (row * 640 + col) <= 161279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161280 && (row * 640 + col) <= 161347) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 161348 && (row * 640 + col) <= 161476) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161477 && (row * 640 + col) <= 161478) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161479 && (row * 640 + col) <= 161483) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 161484 && (row * 640 + col) <= 161486) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 161487 && (row * 640 + col) <= 161489) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 161490 && (row * 640 + col) <= 161491) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 161492 && (row * 640 + col) <= 161493) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 161494 && (row * 640 + col) <= 161498) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 161499 && (row * 640 + col) <= 161499) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 161500 && (row * 640 + col) <= 161503) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 161504 && (row * 640 + col) <= 161506) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 161507 && (row * 640 + col) <= 161508) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 161509 && (row * 640 + col) <= 161512) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 161513 && (row * 640 + col) <= 161514) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161515 && (row * 640 + col) <= 161557) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161558 && (row * 640 + col) <= 161566) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161567 && (row * 640 + col) <= 161575) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161576 && (row * 640 + col) <= 161581) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161582 && (row * 640 + col) <= 161587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161588 && (row * 640 + col) <= 161602) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161603 && (row * 640 + col) <= 161605) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161606 && (row * 640 + col) <= 161617) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161618 && (row * 640 + col) <= 161626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161627 && (row * 640 + col) <= 161632) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161633 && (row * 640 + col) <= 161644) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161645 && (row * 640 + col) <= 161650) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161651 && (row * 640 + col) <= 161653) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161654 && (row * 640 + col) <= 161659) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161660 && (row * 640 + col) <= 161662) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161663 && (row * 640 + col) <= 161677) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161678 && (row * 640 + col) <= 161678) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161679 && (row * 640 + col) <= 161680) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161681 && (row * 640 + col) <= 161686) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161687 && (row * 640 + col) <= 161689) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161690 && (row * 640 + col) <= 161692) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161693 && (row * 640 + col) <= 161695) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161696 && (row * 640 + col) <= 161701) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161702 && (row * 640 + col) <= 161704) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161705 && (row * 640 + col) <= 161716) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161717 && (row * 640 + col) <= 161722) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161723 && (row * 640 + col) <= 161728) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 161729 && (row * 640 + col) <= 161919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161920 && (row * 640 + col) <= 161988) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 161989 && (row * 640 + col) <= 162116) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162117 && (row * 640 + col) <= 162118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162119 && (row * 640 + col) <= 162125) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162126 && (row * 640 + col) <= 162127) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162128 && (row * 640 + col) <= 162129) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162130 && (row * 640 + col) <= 162131) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162132 && (row * 640 + col) <= 162133) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162134 && (row * 640 + col) <= 162135) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162136 && (row * 640 + col) <= 162136) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162137 && (row * 640 + col) <= 162138) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162139 && (row * 640 + col) <= 162139) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162140 && (row * 640 + col) <= 162141) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162142 && (row * 640 + col) <= 162142) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162143 && (row * 640 + col) <= 162144) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162145 && (row * 640 + col) <= 162146) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162147 && (row * 640 + col) <= 162148) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162149 && (row * 640 + col) <= 162152) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162153 && (row * 640 + col) <= 162154) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162155 && (row * 640 + col) <= 162197) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162198 && (row * 640 + col) <= 162206) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162207 && (row * 640 + col) <= 162215) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162216 && (row * 640 + col) <= 162221) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162222 && (row * 640 + col) <= 162227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162228 && (row * 640 + col) <= 162242) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162243 && (row * 640 + col) <= 162245) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162246 && (row * 640 + col) <= 162257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162258 && (row * 640 + col) <= 162266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162267 && (row * 640 + col) <= 162272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162273 && (row * 640 + col) <= 162284) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162285 && (row * 640 + col) <= 162290) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162291 && (row * 640 + col) <= 162293) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162294 && (row * 640 + col) <= 162299) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162300 && (row * 640 + col) <= 162302) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162303 && (row * 640 + col) <= 162317) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162318 && (row * 640 + col) <= 162318) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162319 && (row * 640 + col) <= 162320) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162321 && (row * 640 + col) <= 162326) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162327 && (row * 640 + col) <= 162329) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162330 && (row * 640 + col) <= 162332) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162333 && (row * 640 + col) <= 162335) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162336 && (row * 640 + col) <= 162341) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162342 && (row * 640 + col) <= 162344) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162345 && (row * 640 + col) <= 162356) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162357 && (row * 640 + col) <= 162362) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162363 && (row * 640 + col) <= 162368) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162369 && (row * 640 + col) <= 162559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162560 && (row * 640 + col) <= 162628) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162629 && (row * 640 + col) <= 162756) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162757 && (row * 640 + col) <= 162758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162759 && (row * 640 + col) <= 162765) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162766 && (row * 640 + col) <= 162767) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162768 && (row * 640 + col) <= 162769) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162770 && (row * 640 + col) <= 162771) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162772 && (row * 640 + col) <= 162773) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162774 && (row * 640 + col) <= 162775) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162776 && (row * 640 + col) <= 162776) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162777 && (row * 640 + col) <= 162778) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162779 && (row * 640 + col) <= 162779) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162780 && (row * 640 + col) <= 162781) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162782 && (row * 640 + col) <= 162782) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162783 && (row * 640 + col) <= 162784) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162785 && (row * 640 + col) <= 162786) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162787 && (row * 640 + col) <= 162788) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 162789 && (row * 640 + col) <= 162792) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 162793 && (row * 640 + col) <= 162794) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162795 && (row * 640 + col) <= 162837) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162838 && (row * 640 + col) <= 162846) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162847 && (row * 640 + col) <= 162855) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162856 && (row * 640 + col) <= 162861) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162862 && (row * 640 + col) <= 162867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162868 && (row * 640 + col) <= 162882) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162883 && (row * 640 + col) <= 162885) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162886 && (row * 640 + col) <= 162897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162898 && (row * 640 + col) <= 162906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162907 && (row * 640 + col) <= 162912) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162913 && (row * 640 + col) <= 162924) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162925 && (row * 640 + col) <= 162930) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162931 && (row * 640 + col) <= 162933) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162934 && (row * 640 + col) <= 162939) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162940 && (row * 640 + col) <= 162942) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162943 && (row * 640 + col) <= 162957) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162958 && (row * 640 + col) <= 162958) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162959 && (row * 640 + col) <= 162960) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162961 && (row * 640 + col) <= 162966) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162967 && (row * 640 + col) <= 162969) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162970 && (row * 640 + col) <= 162972) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162973 && (row * 640 + col) <= 162975) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162976 && (row * 640 + col) <= 162981) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162982 && (row * 640 + col) <= 162984) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162985 && (row * 640 + col) <= 162996) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 162997 && (row * 640 + col) <= 163002) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163003 && (row * 640 + col) <= 163008) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163009 && (row * 640 + col) <= 163199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163200 && (row * 640 + col) <= 163279) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 163280 && (row * 640 + col) <= 163396) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163397 && (row * 640 + col) <= 163398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163399 && (row * 640 + col) <= 163402) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163403 && (row * 640 + col) <= 163404) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163405 && (row * 640 + col) <= 163405) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163406 && (row * 640 + col) <= 163407) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163408 && (row * 640 + col) <= 163409) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163410 && (row * 640 + col) <= 163411) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163412 && (row * 640 + col) <= 163413) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163414 && (row * 640 + col) <= 163415) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163416 && (row * 640 + col) <= 163416) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163417 && (row * 640 + col) <= 163418) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163419 && (row * 640 + col) <= 163419) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163420 && (row * 640 + col) <= 163421) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163422 && (row * 640 + col) <= 163422) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163423 && (row * 640 + col) <= 163424) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163425 && (row * 640 + col) <= 163426) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163427 && (row * 640 + col) <= 163428) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 163429 && (row * 640 + col) <= 163432) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 163433 && (row * 640 + col) <= 163434) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163435 && (row * 640 + col) <= 163483) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163484 && (row * 640 + col) <= 163489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163490 && (row * 640 + col) <= 163495) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163496 && (row * 640 + col) <= 163501) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163502 && (row * 640 + col) <= 163507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163508 && (row * 640 + col) <= 163513) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163514 && (row * 640 + col) <= 163516) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163517 && (row * 640 + col) <= 163522) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163523 && (row * 640 + col) <= 163525) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163526 && (row * 640 + col) <= 163531) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163532 && (row * 640 + col) <= 163534) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163535 && (row * 640 + col) <= 163540) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163541 && (row * 640 + col) <= 163546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163547 && (row * 640 + col) <= 163552) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163553 && (row * 640 + col) <= 163564) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163565 && (row * 640 + col) <= 163570) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163571 && (row * 640 + col) <= 163573) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163574 && (row * 640 + col) <= 163579) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163580 && (row * 640 + col) <= 163582) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163583 && (row * 640 + col) <= 163588) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163589 && (row * 640 + col) <= 163591) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163592 && (row * 640 + col) <= 163597) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163598 && (row * 640 + col) <= 163598) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163599 && (row * 640 + col) <= 163600) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 163601 && (row * 640 + col) <= 163606) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163607 && (row * 640 + col) <= 163615) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163616 && (row * 640 + col) <= 163621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163622 && (row * 640 + col) <= 163624) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163625 && (row * 640 + col) <= 163630) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163631 && (row * 640 + col) <= 163642) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163643 && (row * 640 + col) <= 163648) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 163649 && (row * 640 + col) <= 163839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163840 && (row * 640 + col) <= 163919) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 163920 && (row * 640 + col) <= 164036) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164037 && (row * 640 + col) <= 164038) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164039 && (row * 640 + col) <= 164042) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164043 && (row * 640 + col) <= 164047) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 164048 && (row * 640 + col) <= 164049) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164050 && (row * 640 + col) <= 164051) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 164052 && (row * 640 + col) <= 164053) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164054 && (row * 640 + col) <= 164055) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 164056 && (row * 640 + col) <= 164056) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164057 && (row * 640 + col) <= 164058) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 164059 && (row * 640 + col) <= 164059) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164060 && (row * 640 + col) <= 164061) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 164062 && (row * 640 + col) <= 164062) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164063 && (row * 640 + col) <= 164064) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 164065 && (row * 640 + col) <= 164066) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164067 && (row * 640 + col) <= 164068) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 164069 && (row * 640 + col) <= 164072) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164073 && (row * 640 + col) <= 164074) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164075 && (row * 640 + col) <= 164123) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164124 && (row * 640 + col) <= 164129) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164130 && (row * 640 + col) <= 164135) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164136 && (row * 640 + col) <= 164141) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164142 && (row * 640 + col) <= 164147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164148 && (row * 640 + col) <= 164153) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164154 && (row * 640 + col) <= 164156) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164157 && (row * 640 + col) <= 164162) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164163 && (row * 640 + col) <= 164165) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164166 && (row * 640 + col) <= 164171) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164172 && (row * 640 + col) <= 164174) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164175 && (row * 640 + col) <= 164180) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164181 && (row * 640 + col) <= 164186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164187 && (row * 640 + col) <= 164192) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164193 && (row * 640 + col) <= 164204) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164205 && (row * 640 + col) <= 164210) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164211 && (row * 640 + col) <= 164213) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164214 && (row * 640 + col) <= 164219) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164220 && (row * 640 + col) <= 164222) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164223 && (row * 640 + col) <= 164228) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164229 && (row * 640 + col) <= 164231) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164232 && (row * 640 + col) <= 164237) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164238 && (row * 640 + col) <= 164238) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164239 && (row * 640 + col) <= 164240) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164241 && (row * 640 + col) <= 164246) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164247 && (row * 640 + col) <= 164255) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164256 && (row * 640 + col) <= 164261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164262 && (row * 640 + col) <= 164264) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164265 && (row * 640 + col) <= 164270) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164271 && (row * 640 + col) <= 164282) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164283 && (row * 640 + col) <= 164288) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164289 && (row * 640 + col) <= 164479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164480 && (row * 640 + col) <= 164558) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164559 && (row * 640 + col) <= 164676) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164677 && (row * 640 + col) <= 164679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164680 && (row * 640 + col) <= 164711) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 164712 && (row * 640 + col) <= 164714) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164715 && (row * 640 + col) <= 164763) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164764 && (row * 640 + col) <= 164769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164770 && (row * 640 + col) <= 164775) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164776 && (row * 640 + col) <= 164781) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164782 && (row * 640 + col) <= 164787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164788 && (row * 640 + col) <= 164793) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164794 && (row * 640 + col) <= 164796) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164797 && (row * 640 + col) <= 164802) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164803 && (row * 640 + col) <= 164805) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164806 && (row * 640 + col) <= 164811) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164812 && (row * 640 + col) <= 164814) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164815 && (row * 640 + col) <= 164820) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164821 && (row * 640 + col) <= 164826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164827 && (row * 640 + col) <= 164832) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164833 && (row * 640 + col) <= 164844) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164845 && (row * 640 + col) <= 164850) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164851 && (row * 640 + col) <= 164853) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164854 && (row * 640 + col) <= 164859) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164860 && (row * 640 + col) <= 164862) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164863 && (row * 640 + col) <= 164868) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164869 && (row * 640 + col) <= 164871) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164872 && (row * 640 + col) <= 164877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164878 && (row * 640 + col) <= 164878) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164879 && (row * 640 + col) <= 164880) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164881 && (row * 640 + col) <= 164886) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164887 && (row * 640 + col) <= 164895) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164896 && (row * 640 + col) <= 164901) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164902 && (row * 640 + col) <= 164904) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164905 && (row * 640 + col) <= 164910) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164911 && (row * 640 + col) <= 164922) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 164923 && (row * 640 + col) <= 164928) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 164929 && (row * 640 + col) <= 165119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165120 && (row * 640 + col) <= 165182) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165183 && (row * 640 + col) <= 165317) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165318 && (row * 640 + col) <= 165319) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165320 && (row * 640 + col) <= 165351) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 165352 && (row * 640 + col) <= 165353) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165354 && (row * 640 + col) <= 165403) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165404 && (row * 640 + col) <= 165409) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165410 && (row * 640 + col) <= 165415) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165416 && (row * 640 + col) <= 165421) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165422 && (row * 640 + col) <= 165427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165428 && (row * 640 + col) <= 165433) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165434 && (row * 640 + col) <= 165436) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165437 && (row * 640 + col) <= 165442) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165443 && (row * 640 + col) <= 165445) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165446 && (row * 640 + col) <= 165451) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165452 && (row * 640 + col) <= 165454) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165455 && (row * 640 + col) <= 165460) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165461 && (row * 640 + col) <= 165466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165467 && (row * 640 + col) <= 165472) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165473 && (row * 640 + col) <= 165484) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165485 && (row * 640 + col) <= 165490) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165491 && (row * 640 + col) <= 165493) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165494 && (row * 640 + col) <= 165499) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165500 && (row * 640 + col) <= 165502) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165503 && (row * 640 + col) <= 165508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165509 && (row * 640 + col) <= 165511) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165512 && (row * 640 + col) <= 165517) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165518 && (row * 640 + col) <= 165518) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165519 && (row * 640 + col) <= 165520) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 165521 && (row * 640 + col) <= 165526) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165527 && (row * 640 + col) <= 165535) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165536 && (row * 640 + col) <= 165541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165542 && (row * 640 + col) <= 165544) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165545 && (row * 640 + col) <= 165550) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165551 && (row * 640 + col) <= 165572) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165573 && (row * 640 + col) <= 165587) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165588 && (row * 640 + col) <= 165759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165760 && (row * 640 + col) <= 165822) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165823 && (row * 640 + col) <= 165957) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 165958 && (row * 640 + col) <= 165959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165960 && (row * 640 + col) <= 165991) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 165992 && (row * 640 + col) <= 165993) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 165994 && (row * 640 + col) <= 166043) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166044 && (row * 640 + col) <= 166049) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166050 && (row * 640 + col) <= 166055) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166056 && (row * 640 + col) <= 166061) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166062 && (row * 640 + col) <= 166067) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166068 && (row * 640 + col) <= 166073) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166074 && (row * 640 + col) <= 166076) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166077 && (row * 640 + col) <= 166082) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166083 && (row * 640 + col) <= 166085) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166086 && (row * 640 + col) <= 166091) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166092 && (row * 640 + col) <= 166094) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166095 && (row * 640 + col) <= 166100) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166101 && (row * 640 + col) <= 166106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166107 && (row * 640 + col) <= 166112) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166113 && (row * 640 + col) <= 166124) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166125 && (row * 640 + col) <= 166130) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166131 && (row * 640 + col) <= 166133) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166134 && (row * 640 + col) <= 166139) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166140 && (row * 640 + col) <= 166142) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166143 && (row * 640 + col) <= 166148) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166149 && (row * 640 + col) <= 166151) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166152 && (row * 640 + col) <= 166157) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166158 && (row * 640 + col) <= 166158) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166159 && (row * 640 + col) <= 166160) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166161 && (row * 640 + col) <= 166166) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166167 && (row * 640 + col) <= 166175) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166176 && (row * 640 + col) <= 166181) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166182 && (row * 640 + col) <= 166184) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166185 && (row * 640 + col) <= 166190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166191 && (row * 640 + col) <= 166212) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166213 && (row * 640 + col) <= 166227) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166228 && (row * 640 + col) <= 166399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166400 && (row * 640 + col) <= 166440) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166441 && (row * 640 + col) <= 166597) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166598 && (row * 640 + col) <= 166600) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166601 && (row * 640 + col) <= 166630) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 166631 && (row * 640 + col) <= 166633) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166634 && (row * 640 + col) <= 166651) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166652 && (row * 640 + col) <= 166655) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166656 && (row * 640 + col) <= 166683) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166684 && (row * 640 + col) <= 166689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166690 && (row * 640 + col) <= 166695) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166696 && (row * 640 + col) <= 166701) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166702 && (row * 640 + col) <= 166707) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166708 && (row * 640 + col) <= 166713) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166714 && (row * 640 + col) <= 166716) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166717 && (row * 640 + col) <= 166722) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166723 && (row * 640 + col) <= 166725) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166726 && (row * 640 + col) <= 166731) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166732 && (row * 640 + col) <= 166734) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166735 && (row * 640 + col) <= 166740) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166741 && (row * 640 + col) <= 166746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166747 && (row * 640 + col) <= 166752) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166753 && (row * 640 + col) <= 166764) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166765 && (row * 640 + col) <= 166770) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166771 && (row * 640 + col) <= 166773) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166774 && (row * 640 + col) <= 166779) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166780 && (row * 640 + col) <= 166782) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166783 && (row * 640 + col) <= 166788) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166789 && (row * 640 + col) <= 166791) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166792 && (row * 640 + col) <= 166797) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166798 && (row * 640 + col) <= 166798) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166799 && (row * 640 + col) <= 166800) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166801 && (row * 640 + col) <= 166806) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166807 && (row * 640 + col) <= 166815) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166816 && (row * 640 + col) <= 166821) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166822 && (row * 640 + col) <= 166824) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166825 && (row * 640 + col) <= 166830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 166831 && (row * 640 + col) <= 166851) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 166852 && (row * 640 + col) <= 166877) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166878 && (row * 640 + col) <= 167039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167040 && (row * 640 + col) <= 167079) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167080 && (row * 640 + col) <= 167238) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167239 && (row * 640 + col) <= 167240) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167241 && (row * 640 + col) <= 167270) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 167271 && (row * 640 + col) <= 167272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167273 && (row * 640 + col) <= 167291) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167292 && (row * 640 + col) <= 167295) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167296 && (row * 640 + col) <= 167314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167315 && (row * 640 + col) <= 167320) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167321 && (row * 640 + col) <= 167323) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167324 && (row * 640 + col) <= 167329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167330 && (row * 640 + col) <= 167335) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167336 && (row * 640 + col) <= 167341) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167342 && (row * 640 + col) <= 167347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167348 && (row * 640 + col) <= 167353) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167354 && (row * 640 + col) <= 167356) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167357 && (row * 640 + col) <= 167362) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167363 && (row * 640 + col) <= 167365) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167366 && (row * 640 + col) <= 167371) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167372 && (row * 640 + col) <= 167374) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167375 && (row * 640 + col) <= 167380) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167381 && (row * 640 + col) <= 167386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167387 && (row * 640 + col) <= 167392) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167393 && (row * 640 + col) <= 167404) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167405 && (row * 640 + col) <= 167410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167411 && (row * 640 + col) <= 167413) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167414 && (row * 640 + col) <= 167419) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167420 && (row * 640 + col) <= 167422) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167423 && (row * 640 + col) <= 167428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167429 && (row * 640 + col) <= 167431) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167432 && (row * 640 + col) <= 167437) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167438 && (row * 640 + col) <= 167438) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167439 && (row * 640 + col) <= 167440) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167441 && (row * 640 + col) <= 167446) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167447 && (row * 640 + col) <= 167455) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167456 && (row * 640 + col) <= 167461) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167462 && (row * 640 + col) <= 167464) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167465 && (row * 640 + col) <= 167470) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167471 && (row * 640 + col) <= 167473) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167474 && (row * 640 + col) <= 167479) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167480 && (row * 640 + col) <= 167482) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167483 && (row * 640 + col) <= 167488) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167489 && (row * 640 + col) <= 167490) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167491 && (row * 640 + col) <= 167518) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167519 && (row * 640 + col) <= 167679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167680 && (row * 640 + col) <= 167719) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167720 && (row * 640 + col) <= 167878) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167879 && (row * 640 + col) <= 167881) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167882 && (row * 640 + col) <= 167909) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 167910 && (row * 640 + col) <= 167912) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167913 && (row * 640 + col) <= 167931) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167932 && (row * 640 + col) <= 167935) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167936 && (row * 640 + col) <= 167954) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167955 && (row * 640 + col) <= 167960) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167961 && (row * 640 + col) <= 167963) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167964 && (row * 640 + col) <= 167969) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167970 && (row * 640 + col) <= 167975) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167976 && (row * 640 + col) <= 167981) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167982 && (row * 640 + col) <= 167987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167988 && (row * 640 + col) <= 167993) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 167994 && (row * 640 + col) <= 167996) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 167997 && (row * 640 + col) <= 168002) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168003 && (row * 640 + col) <= 168005) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168006 && (row * 640 + col) <= 168011) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168012 && (row * 640 + col) <= 168014) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168015 && (row * 640 + col) <= 168020) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168021 && (row * 640 + col) <= 168026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168027 && (row * 640 + col) <= 168032) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168033 && (row * 640 + col) <= 168044) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168045 && (row * 640 + col) <= 168050) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168051 && (row * 640 + col) <= 168053) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168054 && (row * 640 + col) <= 168059) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168060 && (row * 640 + col) <= 168062) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168063 && (row * 640 + col) <= 168068) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168069 && (row * 640 + col) <= 168071) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168072 && (row * 640 + col) <= 168077) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168078 && (row * 640 + col) <= 168078) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168079 && (row * 640 + col) <= 168080) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 168081 && (row * 640 + col) <= 168086) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168087 && (row * 640 + col) <= 168095) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168096 && (row * 640 + col) <= 168101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168102 && (row * 640 + col) <= 168104) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168105 && (row * 640 + col) <= 168110) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168111 && (row * 640 + col) <= 168113) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168114 && (row * 640 + col) <= 168119) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168120 && (row * 640 + col) <= 168122) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168123 && (row * 640 + col) <= 168128) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168129 && (row * 640 + col) <= 168129) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168130 && (row * 640 + col) <= 168158) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 168159 && (row * 640 + col) <= 168519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168520 && (row * 640 + col) <= 168522) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168523 && (row * 640 + col) <= 168548) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 168549 && (row * 640 + col) <= 168551) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168552 && (row * 640 + col) <= 168571) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168572 && (row * 640 + col) <= 168575) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168576 && (row * 640 + col) <= 168594) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168595 && (row * 640 + col) <= 168600) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168601 && (row * 640 + col) <= 168603) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168604 && (row * 640 + col) <= 168609) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168610 && (row * 640 + col) <= 168615) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168616 && (row * 640 + col) <= 168621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168622 && (row * 640 + col) <= 168627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168628 && (row * 640 + col) <= 168633) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168634 && (row * 640 + col) <= 168636) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168637 && (row * 640 + col) <= 168642) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168643 && (row * 640 + col) <= 168645) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168646 && (row * 640 + col) <= 168651) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168652 && (row * 640 + col) <= 168654) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168655 && (row * 640 + col) <= 168660) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168661 && (row * 640 + col) <= 168666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168667 && (row * 640 + col) <= 168672) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168673 && (row * 640 + col) <= 168684) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168685 && (row * 640 + col) <= 168690) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168691 && (row * 640 + col) <= 168693) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168694 && (row * 640 + col) <= 168699) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168700 && (row * 640 + col) <= 168702) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168703 && (row * 640 + col) <= 168708) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168709 && (row * 640 + col) <= 168711) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168712 && (row * 640 + col) <= 168717) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168718 && (row * 640 + col) <= 168718) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168719 && (row * 640 + col) <= 168720) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 168721 && (row * 640 + col) <= 168726) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168727 && (row * 640 + col) <= 168735) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168736 && (row * 640 + col) <= 168741) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168742 && (row * 640 + col) <= 168744) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168745 && (row * 640 + col) <= 168750) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168751 && (row * 640 + col) <= 168753) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168754 && (row * 640 + col) <= 168759) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168760 && (row * 640 + col) <= 168762) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 168763 && (row * 640 + col) <= 168768) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 168769 && (row * 640 + col) <= 168803) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 168804 && (row * 640 + col) <= 169160) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169161 && (row * 640 + col) <= 169163) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169164 && (row * 640 + col) <= 169187) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 169188 && (row * 640 + col) <= 169190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169191 && (row * 640 + col) <= 169234) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169235 && (row * 640 + col) <= 169249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169250 && (row * 640 + col) <= 169255) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169256 && (row * 640 + col) <= 169261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169262 && (row * 640 + col) <= 169267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169268 && (row * 640 + col) <= 169273) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169274 && (row * 640 + col) <= 169276) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169277 && (row * 640 + col) <= 169282) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169283 && (row * 640 + col) <= 169285) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169286 && (row * 640 + col) <= 169291) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169292 && (row * 640 + col) <= 169294) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169295 && (row * 640 + col) <= 169300) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169301 && (row * 640 + col) <= 169306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169307 && (row * 640 + col) <= 169312) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169313 && (row * 640 + col) <= 169324) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169325 && (row * 640 + col) <= 169339) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169340 && (row * 640 + col) <= 169342) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169343 && (row * 640 + col) <= 169348) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169349 && (row * 640 + col) <= 169351) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169352 && (row * 640 + col) <= 169357) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169358 && (row * 640 + col) <= 169358) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169359 && (row * 640 + col) <= 169360) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 169361 && (row * 640 + col) <= 169366) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169367 && (row * 640 + col) <= 169375) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169376 && (row * 640 + col) <= 169381) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169382 && (row * 640 + col) <= 169384) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169385 && (row * 640 + col) <= 169399) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169400 && (row * 640 + col) <= 169402) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169403 && (row * 640 + col) <= 169408) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169409 && (row * 640 + col) <= 169444) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 169445 && (row * 640 + col) <= 169801) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169802 && (row * 640 + col) <= 169804) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169805 && (row * 640 + col) <= 169826) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 169827 && (row * 640 + col) <= 169829) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169830 && (row * 640 + col) <= 169874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169875 && (row * 640 + col) <= 169889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169890 && (row * 640 + col) <= 169895) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169896 && (row * 640 + col) <= 169901) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169902 && (row * 640 + col) <= 169907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169908 && (row * 640 + col) <= 169913) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169914 && (row * 640 + col) <= 169916) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169917 && (row * 640 + col) <= 169922) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169923 && (row * 640 + col) <= 169925) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169926 && (row * 640 + col) <= 169931) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169932 && (row * 640 + col) <= 169934) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169935 && (row * 640 + col) <= 169940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169941 && (row * 640 + col) <= 169946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169947 && (row * 640 + col) <= 169952) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169953 && (row * 640 + col) <= 169964) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169965 && (row * 640 + col) <= 169979) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169980 && (row * 640 + col) <= 169982) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169983 && (row * 640 + col) <= 169988) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169989 && (row * 640 + col) <= 169991) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169992 && (row * 640 + col) <= 169997) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 169998 && (row * 640 + col) <= 169998) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 169999 && (row * 640 + col) <= 170000) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 170001 && (row * 640 + col) <= 170006) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170007 && (row * 640 + col) <= 170015) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170016 && (row * 640 + col) <= 170021) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170022 && (row * 640 + col) <= 170024) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170025 && (row * 640 + col) <= 170039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170040 && (row * 640 + col) <= 170042) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170043 && (row * 640 + col) <= 170048) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170049 && (row * 640 + col) <= 170084) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 170085 && (row * 640 + col) <= 170442) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170443 && (row * 640 + col) <= 170445) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170446 && (row * 640 + col) <= 170465) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 170466 && (row * 640 + col) <= 170468) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170469 && (row * 640 + col) <= 170514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170515 && (row * 640 + col) <= 170529) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170530 && (row * 640 + col) <= 170535) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170536 && (row * 640 + col) <= 170541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170542 && (row * 640 + col) <= 170547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170548 && (row * 640 + col) <= 170553) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170554 && (row * 640 + col) <= 170556) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170557 && (row * 640 + col) <= 170562) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170563 && (row * 640 + col) <= 170565) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170566 && (row * 640 + col) <= 170571) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170572 && (row * 640 + col) <= 170574) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170575 && (row * 640 + col) <= 170580) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170581 && (row * 640 + col) <= 170586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170587 && (row * 640 + col) <= 170592) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170593 && (row * 640 + col) <= 170604) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170605 && (row * 640 + col) <= 170619) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170620 && (row * 640 + col) <= 170622) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170623 && (row * 640 + col) <= 170628) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170629 && (row * 640 + col) <= 170631) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170632 && (row * 640 + col) <= 170637) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170638 && (row * 640 + col) <= 170640) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 170641 && (row * 640 + col) <= 170646) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170647 && (row * 640 + col) <= 170655) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170656 && (row * 640 + col) <= 170661) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170662 && (row * 640 + col) <= 170664) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170665 && (row * 640 + col) <= 170679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170680 && (row * 640 + col) <= 170682) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 170683 && (row * 640 + col) <= 170688) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 170689 && (row * 640 + col) <= 170726) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 170727 && (row * 640 + col) <= 171083) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 171084 && (row * 640 + col) <= 171086) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 171087 && (row * 640 + col) <= 171104) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 171105 && (row * 640 + col) <= 171107) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 171108 && (row * 640 + col) <= 171272) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 171273 && (row * 640 + col) <= 171286) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171287 && (row * 640 + col) <= 171321) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 171322 && (row * 640 + col) <= 171367) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 171368 && (row * 640 + col) <= 171724) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 171725 && (row * 640 + col) <= 171728) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 171729 && (row * 640 + col) <= 171742) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 171743 && (row * 640 + col) <= 171746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 171747 && (row * 640 + col) <= 171912) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 171913 && (row * 640 + col) <= 171927) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171928 && (row * 640 + col) <= 171961) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 171962 && (row * 640 + col) <= 172007) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 172008 && (row * 640 + col) <= 172365) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 172366 && (row * 640 + col) <= 172371) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 172372 && (row * 640 + col) <= 172379) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 172380 && (row * 640 + col) <= 172385) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 172386 && (row * 640 + col) <= 172552) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 172553 && (row * 640 + col) <= 172567) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 172568 && (row * 640 + col) <= 172598) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 172599 && (row * 640 + col) <= 172647) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 172648 && (row * 640 + col) <= 173007) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 173008 && (row * 640 + col) <= 173023) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 173024 && (row * 640 + col) <= 173192) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 173193 && (row * 640 + col) <= 173206) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173207 && (row * 640 + col) <= 173238) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 173239 && (row * 640 + col) <= 173287) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173288 && (row * 640 + col) <= 173650) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 173651 && (row * 640 + col) <= 173660) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 173661 && (row * 640 + col) <= 173832) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 173833 && (row * 640 + col) <= 173847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173848 && (row * 640 + col) <= 173878) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 173879 && (row * 640 + col) <= 173927) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173928 && (row * 640 + col) <= 174466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 174467 && (row * 640 + col) <= 174492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 174493 && (row * 640 + col) <= 174516) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 174517 && (row * 640 + col) <= 174569) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 174570 && (row * 640 + col) <= 175106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 175107 && (row * 640 + col) <= 175132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 175133 && (row * 640 + col) <= 175155) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 175156 && (row * 640 + col) <= 175210) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 175211 && (row * 640 + col) <= 175746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 175747 && (row * 640 + col) <= 175772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 175773 && (row * 640 + col) <= 175795) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 175796 && (row * 640 + col) <= 175850) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 175851 && (row * 640 + col) <= 176386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 176387 && (row * 640 + col) <= 176412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 176413 && (row * 640 + col) <= 176427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 176428 && (row * 640 + col) <= 176490) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 176491 && (row * 640 + col) <= 177026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 177027 && (row * 640 + col) <= 177052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 177053 && (row * 640 + col) <= 177066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 177067 && (row * 640 + col) <= 177130) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 177131 && (row * 640 + col) <= 177666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 177667 && (row * 640 + col) <= 177692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 177693 && (row * 640 + col) <= 177706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 177707 && (row * 640 + col) <= 177770) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 177771 && (row * 640 + col) <= 178306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 178307 && (row * 640 + col) <= 178332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 178333 && (row * 640 + col) <= 178341) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 178342 && (row * 640 + col) <= 178410) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 178411 && (row * 640 + col) <= 178946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 178947 && (row * 640 + col) <= 178972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 178973 && (row * 640 + col) <= 178981) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 178982 && (row * 640 + col) <= 179050) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 179051 && (row * 640 + col) <= 179586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 179587 && (row * 640 + col) <= 179612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 179613 && (row * 640 + col) <= 179620) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 179621 && (row * 640 + col) <= 179690) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 179691 && (row * 640 + col) <= 180226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 180227 && (row * 640 + col) <= 180252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 180253 && (row * 640 + col) <= 180258) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 180259 && (row * 640 + col) <= 180335) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 180336 && (row * 640 + col) <= 180866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 180867 && (row * 640 + col) <= 180892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 180893 && (row * 640 + col) <= 180898) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 180899 && (row * 640 + col) <= 180976) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 180977 && (row * 640 + col) <= 181506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 181507 && (row * 640 + col) <= 181532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 181533 && (row * 640 + col) <= 181538) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 181539 && (row * 640 + col) <= 181617) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 181618 && (row * 640 + col) <= 182146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 182147 && (row * 640 + col) <= 182172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 182173 && (row * 640 + col) <= 182178) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 182179 && (row * 640 + col) <= 182258) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 182259 && (row * 640 + col) <= 182786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 182787 && (row * 640 + col) <= 182812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 182813 && (row * 640 + col) <= 182818) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 182819 && (row * 640 + col) <= 182898) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 182899 && (row * 640 + col) <= 183426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 183427 && (row * 640 + col) <= 183452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 183453 && (row * 640 + col) <= 183456) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 183457 && (row * 640 + col) <= 183543) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 183544 && (row * 640 + col) <= 184066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 184067 && (row * 640 + col) <= 184092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 184093 && (row * 640 + col) <= 184095) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 184096 && (row * 640 + col) <= 184184) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 184185 && (row * 640 + col) <= 184706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 184707 && (row * 640 + col) <= 184732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 184733 && (row * 640 + col) <= 184735) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 184736 && (row * 640 + col) <= 184824) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 184825 && (row * 640 + col) <= 185346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 185347 && (row * 640 + col) <= 185372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 185373 && (row * 640 + col) <= 185373) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 185374 && (row * 640 + col) <= 185466) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 185467 && (row * 640 + col) <= 185986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 185987 && (row * 640 + col) <= 186012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 186013 && (row * 640 + col) <= 186107) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 186108 && (row * 640 + col) <= 186626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 186627 && (row * 640 + col) <= 186652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 186653 && (row * 640 + col) <= 186747) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 186748 && (row * 640 + col) <= 187266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 187267 && (row * 640 + col) <= 187292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 187293 && (row * 640 + col) <= 187392) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 187393 && (row * 640 + col) <= 187906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 187907 && (row * 640 + col) <= 187932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 187933 && (row * 640 + col) <= 188033) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 188034 && (row * 640 + col) <= 188546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 188547 && (row * 640 + col) <= 188572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 188573 && (row * 640 + col) <= 188672) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 188673 && (row * 640 + col) <= 189186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 189187 && (row * 640 + col) <= 189212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 189213 && (row * 640 + col) <= 189230) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 189231 && (row * 640 + col) <= 189244) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 189245 && (row * 640 + col) <= 189298) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 189299 && (row * 640 + col) <= 189826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 189827 && (row * 640 + col) <= 189852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 189853 && (row * 640 + col) <= 189869) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 189870 && (row * 640 + col) <= 189884) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 189885 && (row * 640 + col) <= 189938) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 189939 && (row * 640 + col) <= 190466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 190467 && (row * 640 + col) <= 190492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 190493 && (row * 640 + col) <= 190493) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 190494 && (row * 640 + col) <= 190509) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 190510 && (row * 640 + col) <= 190524) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 190525 && (row * 640 + col) <= 190528) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 190529 && (row * 640 + col) <= 190530) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 190531 && (row * 640 + col) <= 190542) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 190543 && (row * 640 + col) <= 190544) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 190545 && (row * 640 + col) <= 190553) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 190554 && (row * 640 + col) <= 190557) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 190558 && (row * 640 + col) <= 190578) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 190579 && (row * 640 + col) <= 191106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191107 && (row * 640 + col) <= 191132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 191133 && (row * 640 + col) <= 191141) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191142 && (row * 640 + col) <= 191143) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 191144 && (row * 640 + col) <= 191165) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191166 && (row * 640 + col) <= 191166) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 191167 && (row * 640 + col) <= 191176) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191177 && (row * 640 + col) <= 191178) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 191179 && (row * 640 + col) <= 191187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191188 && (row * 640 + col) <= 191189) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 191190 && (row * 640 + col) <= 191199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191200 && (row * 640 + col) <= 191200) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 191201 && (row * 640 + col) <= 191210) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191211 && (row * 640 + col) <= 191212) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 191213 && (row * 640 + col) <= 191746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 191747 && (row * 640 + col) <= 191772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 191773 && (row * 640 + col) <= 192386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 192387 && (row * 640 + col) <= 192412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 192413 && (row * 640 + col) <= 192812) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 192813 && (row * 640 + col) <= 192828) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 192829 && (row * 640 + col) <= 192986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 192987 && (row * 640 + col) <= 193006) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 193007 && (row * 640 + col) <= 193026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 193027 && (row * 640 + col) <= 193052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 193053 && (row * 640 + col) <= 193446) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 193447 && (row * 640 + col) <= 193472) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 193473 && (row * 640 + col) <= 193626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 193627 && (row * 640 + col) <= 193646) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 193647 && (row * 640 + col) <= 193666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 193667 && (row * 640 + col) <= 193692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 193693 && (row * 640 + col) <= 194082) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 194083 && (row * 640 + col) <= 194093) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 194094 && (row * 640 + col) <= 194107) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 194108 && (row * 640 + col) <= 194114) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 194115 && (row * 640 + col) <= 194266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 194267 && (row * 640 + col) <= 194286) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 194287 && (row * 640 + col) <= 194306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 194307 && (row * 640 + col) <= 194332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 194333 && (row * 640 + col) <= 194718) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 194719 && (row * 640 + col) <= 194727) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 194728 && (row * 640 + col) <= 194751) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 194752 && (row * 640 + col) <= 194757) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 194758 && (row * 640 + col) <= 194906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 194907 && (row * 640 + col) <= 194926) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 194927 && (row * 640 + col) <= 194946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 194947 && (row * 640 + col) <= 194972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 194973 && (row * 640 + col) <= 195356) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 195357 && (row * 640 + col) <= 195363) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 195364 && (row * 640 + col) <= 195393) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 195394 && (row * 640 + col) <= 195400) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 195401 && (row * 640 + col) <= 195546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 195547 && (row * 640 + col) <= 195566) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 195567 && (row * 640 + col) <= 195586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 195587 && (row * 640 + col) <= 195612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 195613 && (row * 640 + col) <= 195995) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 195996 && (row * 640 + col) <= 195999) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 196000 && (row * 640 + col) <= 196036) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 196037 && (row * 640 + col) <= 196043) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 196044 && (row * 640 + col) <= 196186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 196187 && (row * 640 + col) <= 196206) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 196207 && (row * 640 + col) <= 196226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 196227 && (row * 640 + col) <= 196252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 196253 && (row * 640 + col) <= 196477) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 196478 && (row * 640 + col) <= 196479) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 196480 && (row * 640 + col) <= 196634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 196635 && (row * 640 + col) <= 196637) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 196638 && (row * 640 + col) <= 196679) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 196680 && (row * 640 + col) <= 196686) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 196687 && (row * 640 + col) <= 196826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 196827 && (row * 640 + col) <= 196846) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 196847 && (row * 640 + col) <= 196866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 196867 && (row * 640 + col) <= 196892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 196893 && (row * 640 + col) <= 197116) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 197117 && (row * 640 + col) <= 197119) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 197120 && (row * 640 + col) <= 197273) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 197274 && (row * 640 + col) <= 197276) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 197277 && (row * 640 + col) <= 197322) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 197323 && (row * 640 + col) <= 197329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 197330 && (row * 640 + col) <= 197466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 197467 && (row * 640 + col) <= 197486) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 197487 && (row * 640 + col) <= 197506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 197507 && (row * 640 + col) <= 197532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 197533 && (row * 640 + col) <= 197756) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 197757 && (row * 640 + col) <= 197759) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 197760 && (row * 640 + col) <= 197912) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 197913 && (row * 640 + col) <= 197915) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 197916 && (row * 640 + col) <= 197949) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 197950 && (row * 640 + col) <= 197959) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 197960 && (row * 640 + col) <= 197965) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 197966 && (row * 640 + col) <= 197971) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 197972 && (row * 640 + col) <= 198106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 198107 && (row * 640 + col) <= 198126) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 198127 && (row * 640 + col) <= 198147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 198148 && (row * 640 + col) <= 198172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 198173 && (row * 640 + col) <= 198394) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 198395 && (row * 640 + col) <= 198399) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 198400 && (row * 640 + col) <= 198551) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 198552 && (row * 640 + col) <= 198554) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 198555 && (row * 640 + col) <= 198589) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 198590 && (row * 640 + col) <= 198599) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 198600 && (row * 640 + col) <= 198608) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 198609 && (row * 640 + col) <= 198613) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 198614 && (row * 640 + col) <= 198746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 198747 && (row * 640 + col) <= 198766) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 198767 && (row * 640 + col) <= 198787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 198788 && (row * 640 + col) <= 198812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 198813 && (row * 640 + col) <= 199032) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199033 && (row * 640 + col) <= 199039) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199040 && (row * 640 + col) <= 199143) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199144 && (row * 640 + col) <= 199145) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199146 && (row * 640 + col) <= 199149) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199150 && (row * 640 + col) <= 199150) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199151 && (row * 640 + col) <= 199160) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199161 && (row * 640 + col) <= 199162) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199163 && (row * 640 + col) <= 199166) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199167 && (row * 640 + col) <= 199167) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199168 && (row * 640 + col) <= 199171) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199172 && (row * 640 + col) <= 199173) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199174 && (row * 640 + col) <= 199177) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199178 && (row * 640 + col) <= 199179) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199180 && (row * 640 + col) <= 199191) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199192 && (row * 640 + col) <= 199193) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 199194 && (row * 640 + col) <= 199236) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 199237 && (row * 640 + col) <= 199239) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 199240 && (row * 640 + col) <= 199250) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 199251 && (row * 640 + col) <= 199254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 199255 && (row * 640 + col) <= 199386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199387 && (row * 640 + col) <= 199406) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 199407 && (row * 640 + col) <= 199427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199428 && (row * 640 + col) <= 199452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 199453 && (row * 640 + col) <= 199671) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199672 && (row * 640 + col) <= 199679) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199680 && (row * 640 + col) <= 199716) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 199717 && (row * 640 + col) <= 199782) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199783 && (row * 640 + col) <= 199793) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199794 && (row * 640 + col) <= 199799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199800 && (row * 640 + col) <= 199820) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 199821 && (row * 640 + col) <= 199831) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199832 && (row * 640 + col) <= 199833) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 199834 && (row * 640 + col) <= 199875) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 199876 && (row * 640 + col) <= 199878) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 199879 && (row * 640 + col) <= 199892) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 199893 && (row * 640 + col) <= 199896) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 199897 && (row * 640 + col) <= 199920) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199921 && (row * 640 + col) <= 199923) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 199924 && (row * 640 + col) <= 199986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 199987 && (row * 640 + col) <= 200014) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200015 && (row * 640 + col) <= 200026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200027 && (row * 640 + col) <= 200046) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200047 && (row * 640 + col) <= 200066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200067 && (row * 640 + col) <= 200092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200093 && (row * 640 + col) <= 200184) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200185 && (row * 640 + col) <= 200207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200208 && (row * 640 + col) <= 200308) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200309 && (row * 640 + col) <= 200319) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 200320 && (row * 640 + col) <= 200356) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200357 && (row * 640 + col) <= 200421) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200422 && (row * 640 + col) <= 200434) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 200435 && (row * 640 + col) <= 200438) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200439 && (row * 640 + col) <= 200460) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 200461 && (row * 640 + col) <= 200471) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200472 && (row * 640 + col) <= 200473) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 200474 && (row * 640 + col) <= 200515) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 200516 && (row * 640 + col) <= 200517) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 200518 && (row * 640 + col) <= 200533) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 200534 && (row * 640 + col) <= 200537) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 200538 && (row * 640 + col) <= 200560) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200561 && (row * 640 + col) <= 200563) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200564 && (row * 640 + col) <= 200626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200627 && (row * 640 + col) <= 200655) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200656 && (row * 640 + col) <= 200666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200667 && (row * 640 + col) <= 200686) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200687 && (row * 640 + col) <= 200706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200707 && (row * 640 + col) <= 200732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200733 && (row * 640 + col) <= 200824) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200825 && (row * 640 + col) <= 200847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200848 && (row * 640 + col) <= 200947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 200948 && (row * 640 + col) <= 200959) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 200960 && (row * 640 + col) <= 200996) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 200997 && (row * 640 + col) <= 201060) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201061 && (row * 640 + col) <= 201074) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 201075 && (row * 640 + col) <= 201078) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201079 && (row * 640 + col) <= 201101) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 201102 && (row * 640 + col) <= 201111) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201112 && (row * 640 + col) <= 201113) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201114 && (row * 640 + col) <= 201154) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 201155 && (row * 640 + col) <= 201157) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 201158 && (row * 640 + col) <= 201175) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 201176 && (row * 640 + col) <= 201178) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201179 && (row * 640 + col) <= 201200) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201201 && (row * 640 + col) <= 201203) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201204 && (row * 640 + col) <= 201266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201267 && (row * 640 + col) <= 201295) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201296 && (row * 640 + col) <= 201306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201307 && (row * 640 + col) <= 201326) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201327 && (row * 640 + col) <= 201346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201347 && (row * 640 + col) <= 201372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201373 && (row * 640 + col) <= 201464) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201465 && (row * 640 + col) <= 201487) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201488 && (row * 640 + col) <= 201587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201588 && (row * 640 + col) <= 201599) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 201600 && (row * 640 + col) <= 201636) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201637 && (row * 640 + col) <= 201696) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201697 && (row * 640 + col) <= 201743) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 201744 && (row * 640 + col) <= 201751) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201752 && (row * 640 + col) <= 201754) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201755 && (row * 640 + col) <= 201794) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 201795 && (row * 640 + col) <= 201796) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 201797 && (row * 640 + col) <= 201816) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 201817 && (row * 640 + col) <= 201820) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201821 && (row * 640 + col) <= 201823) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201824 && (row * 640 + col) <= 201840) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201841 && (row * 640 + col) <= 201843) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201844 && (row * 640 + col) <= 201874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201875 && (row * 640 + col) <= 201886) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201887 && (row * 640 + col) <= 201889) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201890 && (row * 640 + col) <= 201895) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201896 && (row * 640 + col) <= 201901) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201902 && (row * 640 + col) <= 201907) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201908 && (row * 640 + col) <= 201910) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201911 && (row * 640 + col) <= 201925) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201926 && (row * 640 + col) <= 201928) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201929 && (row * 640 + col) <= 201940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201941 && (row * 640 + col) <= 201943) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201944 && (row * 640 + col) <= 201958) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201959 && (row * 640 + col) <= 201961) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201962 && (row * 640 + col) <= 201967) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201968 && (row * 640 + col) <= 201970) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201971 && (row * 640 + col) <= 201976) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201977 && (row * 640 + col) <= 201979) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 201980 && (row * 640 + col) <= 201994) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 201995 && (row * 640 + col) <= 201997) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 201998 && (row * 640 + col) <= 202009) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202010 && (row * 640 + col) <= 202012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202013 && (row * 640 + col) <= 202024) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202025 && (row * 640 + col) <= 202027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202028 && (row * 640 + col) <= 202042) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202043 && (row * 640 + col) <= 202045) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202046 && (row * 640 + col) <= 202051) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202052 && (row * 640 + col) <= 202057) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202058 && (row * 640 + col) <= 202063) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202064 && (row * 640 + col) <= 202066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202067 && (row * 640 + col) <= 202081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202082 && (row * 640 + col) <= 202104) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202105 && (row * 640 + col) <= 202127) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202128 && (row * 640 + col) <= 202221) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202222 && (row * 640 + col) <= 202239) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 202240 && (row * 640 + col) <= 202276) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202277 && (row * 640 + col) <= 202336) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202337 && (row * 640 + col) <= 202383) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 202384 && (row * 640 + col) <= 202392) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202393 && (row * 640 + col) <= 202394) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202395 && (row * 640 + col) <= 202433) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 202434 && (row * 640 + col) <= 202436) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 202437 && (row * 640 + col) <= 202458) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 202459 && (row * 640 + col) <= 202461) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202462 && (row * 640 + col) <= 202463) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202464 && (row * 640 + col) <= 202480) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202481 && (row * 640 + col) <= 202483) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202484 && (row * 640 + col) <= 202514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202515 && (row * 640 + col) <= 202526) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202527 && (row * 640 + col) <= 202529) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202530 && (row * 640 + col) <= 202535) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202536 && (row * 640 + col) <= 202541) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202542 && (row * 640 + col) <= 202547) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202548 && (row * 640 + col) <= 202550) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202551 && (row * 640 + col) <= 202565) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202566 && (row * 640 + col) <= 202568) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202569 && (row * 640 + col) <= 202580) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202581 && (row * 640 + col) <= 202583) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202584 && (row * 640 + col) <= 202598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202599 && (row * 640 + col) <= 202601) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202602 && (row * 640 + col) <= 202607) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202608 && (row * 640 + col) <= 202610) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202611 && (row * 640 + col) <= 202616) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202617 && (row * 640 + col) <= 202619) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202620 && (row * 640 + col) <= 202634) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202635 && (row * 640 + col) <= 202637) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202638 && (row * 640 + col) <= 202649) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202650 && (row * 640 + col) <= 202652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202653 && (row * 640 + col) <= 202664) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202665 && (row * 640 + col) <= 202667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202668 && (row * 640 + col) <= 202682) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202683 && (row * 640 + col) <= 202685) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202686 && (row * 640 + col) <= 202691) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202692 && (row * 640 + col) <= 202697) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202698 && (row * 640 + col) <= 202703) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202704 && (row * 640 + col) <= 202706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202707 && (row * 640 + col) <= 202721) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 202722 && (row * 640 + col) <= 202744) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202745 && (row * 640 + col) <= 202767) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202768 && (row * 640 + col) <= 202860) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202861 && (row * 640 + col) <= 202879) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 202880 && (row * 640 + col) <= 202916) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 202917 && (row * 640 + col) <= 202974) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 202975 && (row * 640 + col) <= 203024) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 203025 && (row * 640 + col) <= 203033) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203034 && (row * 640 + col) <= 203035) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203036 && (row * 640 + col) <= 203072) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 203073 && (row * 640 + col) <= 203075) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 203076 && (row * 640 + col) <= 203099) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 203100 && (row * 640 + col) <= 203102) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203103 && (row * 640 + col) <= 203103) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203104 && (row * 640 + col) <= 203120) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203121 && (row * 640 + col) <= 203123) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203124 && (row * 640 + col) <= 203154) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203155 && (row * 640 + col) <= 203166) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203167 && (row * 640 + col) <= 203169) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203170 && (row * 640 + col) <= 203175) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203176 && (row * 640 + col) <= 203181) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203182 && (row * 640 + col) <= 203187) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203188 && (row * 640 + col) <= 203190) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203191 && (row * 640 + col) <= 203205) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203206 && (row * 640 + col) <= 203208) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203209 && (row * 640 + col) <= 203220) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203221 && (row * 640 + col) <= 203223) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203224 && (row * 640 + col) <= 203238) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203239 && (row * 640 + col) <= 203241) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203242 && (row * 640 + col) <= 203247) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203248 && (row * 640 + col) <= 203250) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203251 && (row * 640 + col) <= 203256) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203257 && (row * 640 + col) <= 203259) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203260 && (row * 640 + col) <= 203274) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203275 && (row * 640 + col) <= 203277) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203278 && (row * 640 + col) <= 203289) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203290 && (row * 640 + col) <= 203292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203293 && (row * 640 + col) <= 203304) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203305 && (row * 640 + col) <= 203307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203308 && (row * 640 + col) <= 203322) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203323 && (row * 640 + col) <= 203325) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203326 && (row * 640 + col) <= 203331) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203332 && (row * 640 + col) <= 203337) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203338 && (row * 640 + col) <= 203343) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203344 && (row * 640 + col) <= 203346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203347 && (row * 640 + col) <= 203361) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203362 && (row * 640 + col) <= 203384) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203385 && (row * 640 + col) <= 203407) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203408 && (row * 640 + col) <= 203490) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203491 && (row * 640 + col) <= 203496) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 203497 && (row * 640 + col) <= 203499) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203500 && (row * 640 + col) <= 203519) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 203520 && (row * 640 + col) <= 203556) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203557 && (row * 640 + col) <= 203613) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203614 && (row * 640 + col) <= 203663) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 203664 && (row * 640 + col) <= 203673) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203674 && (row * 640 + col) <= 203676) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203677 && (row * 640 + col) <= 203712) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 203713 && (row * 640 + col) <= 203714) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 203715 && (row * 640 + col) <= 203740) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 203741 && (row * 640 + col) <= 203743) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203744 && (row * 640 + col) <= 203757) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203758 && (row * 640 + col) <= 203765) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203766 && (row * 640 + col) <= 203771) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203772 && (row * 640 + col) <= 203775) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203776 && (row * 640 + col) <= 203797) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203798 && (row * 640 + col) <= 203803) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203804 && (row * 640 + col) <= 203809) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203810 && (row * 640 + col) <= 203818) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203819 && (row * 640 + col) <= 203821) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203822 && (row * 640 + col) <= 203827) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203828 && (row * 640 + col) <= 203830) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203831 && (row * 640 + col) <= 203836) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203837 && (row * 640 + col) <= 203839) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203840 && (row * 640 + col) <= 203845) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203846 && (row * 640 + col) <= 203851) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203852 && (row * 640 + col) <= 203857) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203858 && (row * 640 + col) <= 203863) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203864 && (row * 640 + col) <= 203869) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203870 && (row * 640 + col) <= 203872) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203873 && (row * 640 + col) <= 203878) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203879 && (row * 640 + col) <= 203881) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203882 && (row * 640 + col) <= 203887) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203888 && (row * 640 + col) <= 203890) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203891 && (row * 640 + col) <= 203896) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203897 && (row * 640 + col) <= 203899) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203900 && (row * 640 + col) <= 203905) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203906 && (row * 640 + col) <= 203907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203908 && (row * 640 + col) <= 203908) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203909 && (row * 640 + col) <= 203914) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203915 && (row * 640 + col) <= 203920) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203921 && (row * 640 + col) <= 203926) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203927 && (row * 640 + col) <= 203932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 203933 && (row * 640 + col) <= 203935) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203936 && (row * 640 + col) <= 203941) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203942 && (row * 640 + col) <= 203947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203948 && (row * 640 + col) <= 203953) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203954 && (row * 640 + col) <= 203956) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203957 && (row * 640 + col) <= 203962) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203963 && (row * 640 + col) <= 203965) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203966 && (row * 640 + col) <= 203974) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203975 && (row * 640 + col) <= 203977) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203978 && (row * 640 + col) <= 203983) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203984 && (row * 640 + col) <= 203986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203987 && (row * 640 + col) <= 203992) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 203993 && (row * 640 + col) <= 203995) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 203996 && (row * 640 + col) <= 204001) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204002 && (row * 640 + col) <= 204018) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204019 && (row * 640 + col) <= 204024) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204025 && (row * 640 + col) <= 204047) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204048 && (row * 640 + col) <= 204129) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204130 && (row * 640 + col) <= 204159) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 204160 && (row * 640 + col) <= 204196) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204197 && (row * 640 + col) <= 204252) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204253 && (row * 640 + col) <= 204303) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 204304 && (row * 640 + col) <= 204314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204315 && (row * 640 + col) <= 204319) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204320 && (row * 640 + col) <= 204351) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 204352 && (row * 640 + col) <= 204354) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 204355 && (row * 640 + col) <= 204381) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 204382 && (row * 640 + col) <= 204384) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204385 && (row * 640 + col) <= 204397) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204398 && (row * 640 + col) <= 204406) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204407 && (row * 640 + col) <= 204411) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204412 && (row * 640 + col) <= 204415) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204416 && (row * 640 + col) <= 204437) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204438 && (row * 640 + col) <= 204443) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204444 && (row * 640 + col) <= 204449) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204450 && (row * 640 + col) <= 204458) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204459 && (row * 640 + col) <= 204461) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204462 && (row * 640 + col) <= 204467) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204468 && (row * 640 + col) <= 204470) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204471 && (row * 640 + col) <= 204476) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204477 && (row * 640 + col) <= 204479) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204480 && (row * 640 + col) <= 204485) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204486 && (row * 640 + col) <= 204491) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204492 && (row * 640 + col) <= 204497) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204498 && (row * 640 + col) <= 204503) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204504 && (row * 640 + col) <= 204509) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204510 && (row * 640 + col) <= 204512) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204513 && (row * 640 + col) <= 204518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204519 && (row * 640 + col) <= 204521) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204522 && (row * 640 + col) <= 204527) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204528 && (row * 640 + col) <= 204530) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204531 && (row * 640 + col) <= 204536) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204537 && (row * 640 + col) <= 204539) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204540 && (row * 640 + col) <= 204545) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204546 && (row * 640 + col) <= 204547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204548 && (row * 640 + col) <= 204548) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204549 && (row * 640 + col) <= 204554) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204555 && (row * 640 + col) <= 204560) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204561 && (row * 640 + col) <= 204566) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204567 && (row * 640 + col) <= 204572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204573 && (row * 640 + col) <= 204575) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204576 && (row * 640 + col) <= 204581) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204582 && (row * 640 + col) <= 204587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204588 && (row * 640 + col) <= 204593) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204594 && (row * 640 + col) <= 204596) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204597 && (row * 640 + col) <= 204602) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204603 && (row * 640 + col) <= 204605) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204606 && (row * 640 + col) <= 204614) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204615 && (row * 640 + col) <= 204617) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204618 && (row * 640 + col) <= 204623) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204624 && (row * 640 + col) <= 204626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204627 && (row * 640 + col) <= 204632) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204633 && (row * 640 + col) <= 204635) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204636 && (row * 640 + col) <= 204641) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204642 && (row * 640 + col) <= 204658) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204659 && (row * 640 + col) <= 204664) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204665 && (row * 640 + col) <= 204687) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204688 && (row * 640 + col) <= 204769) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204770 && (row * 640 + col) <= 204799) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 204800 && (row * 640 + col) <= 204836) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 204837 && (row * 640 + col) <= 204890) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204891 && (row * 640 + col) <= 204944) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 204945 && (row * 640 + col) <= 204955) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 204956 && (row * 640 + col) <= 204965) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 204966 && (row * 640 + col) <= 204991) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 204992 && (row * 640 + col) <= 204993) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 204994 && (row * 640 + col) <= 205022) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 205023 && (row * 640 + col) <= 205025) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205026 && (row * 640 + col) <= 205037) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205038 && (row * 640 + col) <= 205046) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205047 && (row * 640 + col) <= 205051) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205052 && (row * 640 + col) <= 205055) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205056 && (row * 640 + col) <= 205077) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205078 && (row * 640 + col) <= 205083) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205084 && (row * 640 + col) <= 205089) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205090 && (row * 640 + col) <= 205098) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205099 && (row * 640 + col) <= 205101) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205102 && (row * 640 + col) <= 205107) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205108 && (row * 640 + col) <= 205110) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205111 && (row * 640 + col) <= 205116) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205117 && (row * 640 + col) <= 205119) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205120 && (row * 640 + col) <= 205125) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205126 && (row * 640 + col) <= 205131) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205132 && (row * 640 + col) <= 205137) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205138 && (row * 640 + col) <= 205143) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205144 && (row * 640 + col) <= 205149) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205150 && (row * 640 + col) <= 205152) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205153 && (row * 640 + col) <= 205158) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205159 && (row * 640 + col) <= 205161) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205162 && (row * 640 + col) <= 205167) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205168 && (row * 640 + col) <= 205170) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205171 && (row * 640 + col) <= 205176) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205177 && (row * 640 + col) <= 205179) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205180 && (row * 640 + col) <= 205185) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205186 && (row * 640 + col) <= 205187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205188 && (row * 640 + col) <= 205188) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205189 && (row * 640 + col) <= 205194) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205195 && (row * 640 + col) <= 205200) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205201 && (row * 640 + col) <= 205206) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205207 && (row * 640 + col) <= 205212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205213 && (row * 640 + col) <= 205215) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205216 && (row * 640 + col) <= 205221) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205222 && (row * 640 + col) <= 205227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205228 && (row * 640 + col) <= 205233) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205234 && (row * 640 + col) <= 205236) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205237 && (row * 640 + col) <= 205242) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205243 && (row * 640 + col) <= 205245) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205246 && (row * 640 + col) <= 205254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205255 && (row * 640 + col) <= 205257) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205258 && (row * 640 + col) <= 205263) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205264 && (row * 640 + col) <= 205266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205267 && (row * 640 + col) <= 205272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205273 && (row * 640 + col) <= 205275) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205276 && (row * 640 + col) <= 205281) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205282 && (row * 640 + col) <= 205298) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205299 && (row * 640 + col) <= 205304) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205305 && (row * 640 + col) <= 205327) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205328 && (row * 640 + col) <= 205402) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205403 && (row * 640 + col) <= 205439) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 205440 && (row * 640 + col) <= 205476) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205477 && (row * 640 + col) <= 205530) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205531 && (row * 640 + col) <= 205583) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 205584 && (row * 640 + col) <= 205598) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205599 && (row * 640 + col) <= 205610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205611 && (row * 640 + col) <= 205630) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 205631 && (row * 640 + col) <= 205633) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 205634 && (row * 640 + col) <= 205663) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 205664 && (row * 640 + col) <= 205666) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205667 && (row * 640 + col) <= 205677) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205678 && (row * 640 + col) <= 205686) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205687 && (row * 640 + col) <= 205691) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205692 && (row * 640 + col) <= 205695) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205696 && (row * 640 + col) <= 205709) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205710 && (row * 640 + col) <= 205717) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205718 && (row * 640 + col) <= 205723) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205724 && (row * 640 + col) <= 205729) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205730 && (row * 640 + col) <= 205747) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205748 && (row * 640 + col) <= 205750) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205751 && (row * 640 + col) <= 205756) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205757 && (row * 640 + col) <= 205771) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205772 && (row * 640 + col) <= 205777) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205778 && (row * 640 + col) <= 205783) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205784 && (row * 640 + col) <= 205789) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205790 && (row * 640 + col) <= 205792) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205793 && (row * 640 + col) <= 205798) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205799 && (row * 640 + col) <= 205801) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205802 && (row * 640 + col) <= 205807) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205808 && (row * 640 + col) <= 205810) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205811 && (row * 640 + col) <= 205816) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205817 && (row * 640 + col) <= 205819) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205820 && (row * 640 + col) <= 205825) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205826 && (row * 640 + col) <= 205827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205828 && (row * 640 + col) <= 205840) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205841 && (row * 640 + col) <= 205846) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205847 && (row * 640 + col) <= 205852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205853 && (row * 640 + col) <= 205855) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205856 && (row * 640 + col) <= 205861) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205862 && (row * 640 + col) <= 205867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205868 && (row * 640 + col) <= 205873) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205874 && (row * 640 + col) <= 205876) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205877 && (row * 640 + col) <= 205882) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205883 && (row * 640 + col) <= 205885) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205886 && (row * 640 + col) <= 205903) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205904 && (row * 640 + col) <= 205906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205907 && (row * 640 + col) <= 205912) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 205913 && (row * 640 + col) <= 205921) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205922 && (row * 640 + col) <= 205938) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205939 && (row * 640 + col) <= 205944) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 205945 && (row * 640 + col) <= 205967) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 205968 && (row * 640 + col) <= 206041) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206042 && (row * 640 + col) <= 206079) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 206080 && (row * 640 + col) <= 206116) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206117 && (row * 640 + col) <= 206169) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206170 && (row * 640 + col) <= 206223) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 206224 && (row * 640 + col) <= 206244) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206245 && (row * 640 + col) <= 206254) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206255 && (row * 640 + col) <= 206269) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 206270 && (row * 640 + col) <= 206272) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 206273 && (row * 640 + col) <= 206304) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 206305 && (row * 640 + col) <= 206307) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206308 && (row * 640 + col) <= 206317) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206318 && (row * 640 + col) <= 206326) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206327 && (row * 640 + col) <= 206349) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206350 && (row * 640 + col) <= 206357) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206358 && (row * 640 + col) <= 206363) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206364 && (row * 640 + col) <= 206369) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206370 && (row * 640 + col) <= 206387) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206388 && (row * 640 + col) <= 206390) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206391 && (row * 640 + col) <= 206396) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206397 && (row * 640 + col) <= 206411) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206412 && (row * 640 + col) <= 206417) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206418 && (row * 640 + col) <= 206423) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206424 && (row * 640 + col) <= 206429) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206430 && (row * 640 + col) <= 206432) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206433 && (row * 640 + col) <= 206438) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206439 && (row * 640 + col) <= 206441) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206442 && (row * 640 + col) <= 206447) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206448 && (row * 640 + col) <= 206450) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206451 && (row * 640 + col) <= 206456) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206457 && (row * 640 + col) <= 206459) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206460 && (row * 640 + col) <= 206465) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206466 && (row * 640 + col) <= 206467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206468 && (row * 640 + col) <= 206480) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206481 && (row * 640 + col) <= 206486) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206487 && (row * 640 + col) <= 206492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206493 && (row * 640 + col) <= 206495) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206496 && (row * 640 + col) <= 206501) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206502 && (row * 640 + col) <= 206507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206508 && (row * 640 + col) <= 206513) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206514 && (row * 640 + col) <= 206516) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206517 && (row * 640 + col) <= 206522) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206523 && (row * 640 + col) <= 206525) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206526 && (row * 640 + col) <= 206543) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206544 && (row * 640 + col) <= 206546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206547 && (row * 640 + col) <= 206552) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206553 && (row * 640 + col) <= 206561) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206562 && (row * 640 + col) <= 206578) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206579 && (row * 640 + col) <= 206584) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206585 && (row * 640 + col) <= 206607) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206608 && (row * 640 + col) <= 206678) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206679 && (row * 640 + col) <= 206679) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 206680 && (row * 640 + col) <= 206680) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206681 && (row * 640 + col) <= 206719) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 206720 && (row * 640 + col) <= 206756) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206757 && (row * 640 + col) <= 206807) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206808 && (row * 640 + col) <= 206863) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 206864 && (row * 640 + col) <= 206889) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206890 && (row * 640 + col) <= 206900) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206901 && (row * 640 + col) <= 206909) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 206910 && (row * 640 + col) <= 206919) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 206920 && (row * 640 + col) <= 206945) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 206946 && (row * 640 + col) <= 206948) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 206949 && (row * 640 + col) <= 206957) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206958 && (row * 640 + col) <= 206966) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206967 && (row * 640 + col) <= 206989) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 206990 && (row * 640 + col) <= 206997) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 206998 && (row * 640 + col) <= 207003) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207004 && (row * 640 + col) <= 207009) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207010 && (row * 640 + col) <= 207027) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207028 && (row * 640 + col) <= 207030) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207031 && (row * 640 + col) <= 207036) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207037 && (row * 640 + col) <= 207051) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207052 && (row * 640 + col) <= 207057) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207058 && (row * 640 + col) <= 207063) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207064 && (row * 640 + col) <= 207069) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207070 && (row * 640 + col) <= 207072) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207073 && (row * 640 + col) <= 207078) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207079 && (row * 640 + col) <= 207081) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207082 && (row * 640 + col) <= 207087) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207088 && (row * 640 + col) <= 207090) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207091 && (row * 640 + col) <= 207096) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207097 && (row * 640 + col) <= 207099) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207100 && (row * 640 + col) <= 207105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207106 && (row * 640 + col) <= 207107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207108 && (row * 640 + col) <= 207120) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207121 && (row * 640 + col) <= 207126) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207127 && (row * 640 + col) <= 207132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207133 && (row * 640 + col) <= 207135) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207136 && (row * 640 + col) <= 207141) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207142 && (row * 640 + col) <= 207147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207148 && (row * 640 + col) <= 207153) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207154 && (row * 640 + col) <= 207156) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207157 && (row * 640 + col) <= 207162) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207163 && (row * 640 + col) <= 207165) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207166 && (row * 640 + col) <= 207183) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207184 && (row * 640 + col) <= 207186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207187 && (row * 640 + col) <= 207192) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207193 && (row * 640 + col) <= 207201) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207202 && (row * 640 + col) <= 207218) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207219 && (row * 640 + col) <= 207224) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207225 && (row * 640 + col) <= 207247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207248 && (row * 640 + col) <= 207313) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207314 && (row * 640 + col) <= 207359) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 207360 && (row * 640 + col) <= 207396) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207397 && (row * 640 + col) <= 207447) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207448 && (row * 640 + col) <= 207503) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 207504 && (row * 640 + col) <= 207531) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207532 && (row * 640 + col) <= 207533) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207534 && (row * 640 + col) <= 207544) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207545 && (row * 640 + col) <= 207549) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 207550 && (row * 640 + col) <= 207559) color_data <= 12'b010000011001; else
        if ((row * 640 + col) >= 207560 && (row * 640 + col) <= 207586) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 207587 && (row * 640 + col) <= 207589) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207590 && (row * 640 + col) <= 207595) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207596 && (row * 640 + col) <= 207609) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207610 && (row * 640 + col) <= 207629) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207630 && (row * 640 + col) <= 207637) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207638 && (row * 640 + col) <= 207643) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207644 && (row * 640 + col) <= 207649) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207650 && (row * 640 + col) <= 207655) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207656 && (row * 640 + col) <= 207658) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207659 && (row * 640 + col) <= 207667) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207668 && (row * 640 + col) <= 207673) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207674 && (row * 640 + col) <= 207682) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207683 && (row * 640 + col) <= 207691) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207692 && (row * 640 + col) <= 207697) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207698 && (row * 640 + col) <= 207703) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207704 && (row * 640 + col) <= 207715) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207716 && (row * 640 + col) <= 207721) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207722 && (row * 640 + col) <= 207727) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207728 && (row * 640 + col) <= 207730) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207731 && (row * 640 + col) <= 207736) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207737 && (row * 640 + col) <= 207739) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207740 && (row * 640 + col) <= 207745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207746 && (row * 640 + col) <= 207747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207748 && (row * 640 + col) <= 207760) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207761 && (row * 640 + col) <= 207766) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207767 && (row * 640 + col) <= 207772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207773 && (row * 640 + col) <= 207775) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207776 && (row * 640 + col) <= 207781) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207782 && (row * 640 + col) <= 207787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207788 && (row * 640 + col) <= 207793) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207794 && (row * 640 + col) <= 207796) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207797 && (row * 640 + col) <= 207802) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207803 && (row * 640 + col) <= 207805) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207806 && (row * 640 + col) <= 207811) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207812 && (row * 640 + col) <= 207814) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207815 && (row * 640 + col) <= 207823) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207824 && (row * 640 + col) <= 207829) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207830 && (row * 640 + col) <= 207838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207839 && (row * 640 + col) <= 207841) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207842 && (row * 640 + col) <= 207858) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207859 && (row * 640 + col) <= 207864) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207865 && (row * 640 + col) <= 207887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 207888 && (row * 640 + col) <= 207952) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 207953 && (row * 640 + col) <= 207999) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 208000 && (row * 640 + col) <= 208036) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208037 && (row * 640 + col) <= 208087) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208088 && (row * 640 + col) <= 208144) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 208145 && (row * 640 + col) <= 208171) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208172 && (row * 640 + col) <= 208179) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208180 && (row * 640 + col) <= 208187) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208188 && (row * 640 + col) <= 208227) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 208228 && (row * 640 + col) <= 208230) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208231 && (row * 640 + col) <= 208235) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208236 && (row * 640 + col) <= 208249) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208250 && (row * 640 + col) <= 208269) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208270 && (row * 640 + col) <= 208277) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208278 && (row * 640 + col) <= 208283) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208284 && (row * 640 + col) <= 208289) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208290 && (row * 640 + col) <= 208295) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208296 && (row * 640 + col) <= 208298) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208299 && (row * 640 + col) <= 208307) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208308 && (row * 640 + col) <= 208313) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208314 && (row * 640 + col) <= 208322) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208323 && (row * 640 + col) <= 208331) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208332 && (row * 640 + col) <= 208337) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208338 && (row * 640 + col) <= 208343) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208344 && (row * 640 + col) <= 208355) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208356 && (row * 640 + col) <= 208361) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208362 && (row * 640 + col) <= 208367) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208368 && (row * 640 + col) <= 208370) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208371 && (row * 640 + col) <= 208376) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208377 && (row * 640 + col) <= 208379) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208380 && (row * 640 + col) <= 208385) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208386 && (row * 640 + col) <= 208387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208388 && (row * 640 + col) <= 208400) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208401 && (row * 640 + col) <= 208406) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208407 && (row * 640 + col) <= 208412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208413 && (row * 640 + col) <= 208415) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208416 && (row * 640 + col) <= 208421) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208422 && (row * 640 + col) <= 208427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208428 && (row * 640 + col) <= 208433) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208434 && (row * 640 + col) <= 208436) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208437 && (row * 640 + col) <= 208442) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208443 && (row * 640 + col) <= 208445) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208446 && (row * 640 + col) <= 208451) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208452 && (row * 640 + col) <= 208454) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208455 && (row * 640 + col) <= 208463) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208464 && (row * 640 + col) <= 208469) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208470 && (row * 640 + col) <= 208478) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208479 && (row * 640 + col) <= 208481) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208482 && (row * 640 + col) <= 208498) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208499 && (row * 640 + col) <= 208504) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208505 && (row * 640 + col) <= 208527) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208528 && (row * 640 + col) <= 208592) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208593 && (row * 640 + col) <= 208639) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 208640 && (row * 640 + col) <= 208676) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208677 && (row * 640 + col) <= 208727) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208728 && (row * 640 + col) <= 208785) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 208786 && (row * 640 + col) <= 208811) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208812 && (row * 640 + col) <= 208823) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208824 && (row * 640 + col) <= 208830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208831 && (row * 640 + col) <= 208868) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 208869 && (row * 640 + col) <= 208871) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208872 && (row * 640 + col) <= 208875) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208876 && (row * 640 + col) <= 208888) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208889 && (row * 640 + col) <= 208909) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208910 && (row * 640 + col) <= 208917) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208918 && (row * 640 + col) <= 208923) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208924 && (row * 640 + col) <= 208929) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208930 && (row * 640 + col) <= 208935) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208936 && (row * 640 + col) <= 208938) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208939 && (row * 640 + col) <= 208947) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208948 && (row * 640 + col) <= 208953) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208954 && (row * 640 + col) <= 208962) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208963 && (row * 640 + col) <= 208971) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 208972 && (row * 640 + col) <= 208977) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208978 && (row * 640 + col) <= 208983) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 208984 && (row * 640 + col) <= 208995) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208996 && (row * 640 + col) <= 209001) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209002 && (row * 640 + col) <= 209007) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209008 && (row * 640 + col) <= 209010) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209011 && (row * 640 + col) <= 209016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209017 && (row * 640 + col) <= 209019) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209020 && (row * 640 + col) <= 209025) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209026 && (row * 640 + col) <= 209027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209028 && (row * 640 + col) <= 209040) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209041 && (row * 640 + col) <= 209046) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209047 && (row * 640 + col) <= 209052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209053 && (row * 640 + col) <= 209055) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209056 && (row * 640 + col) <= 209061) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209062 && (row * 640 + col) <= 209067) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209068 && (row * 640 + col) <= 209073) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209074 && (row * 640 + col) <= 209076) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209077 && (row * 640 + col) <= 209082) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209083 && (row * 640 + col) <= 209085) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209086 && (row * 640 + col) <= 209091) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209092 && (row * 640 + col) <= 209094) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209095 && (row * 640 + col) <= 209103) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209104 && (row * 640 + col) <= 209109) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209110 && (row * 640 + col) <= 209118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209119 && (row * 640 + col) <= 209121) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209122 && (row * 640 + col) <= 209138) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209139 && (row * 640 + col) <= 209144) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209145 && (row * 640 + col) <= 209167) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209168 && (row * 640 + col) <= 209230) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209231 && (row * 640 + col) <= 209279) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 209280 && (row * 640 + col) <= 209316) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209317 && (row * 640 + col) <= 209367) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209368 && (row * 640 + col) <= 209426) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 209427 && (row * 640 + col) <= 209451) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209452 && (row * 640 + col) <= 209466) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209467 && (row * 640 + col) <= 209473) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209474 && (row * 640 + col) <= 209509) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 209510 && (row * 640 + col) <= 209511) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209512 && (row * 640 + col) <= 209515) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209516 && (row * 640 + col) <= 209528) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209529 && (row * 640 + col) <= 209549) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209550 && (row * 640 + col) <= 209557) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209558 && (row * 640 + col) <= 209563) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209564 && (row * 640 + col) <= 209569) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209570 && (row * 640 + col) <= 209575) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209576 && (row * 640 + col) <= 209581) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209582 && (row * 640 + col) <= 209587) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209588 && (row * 640 + col) <= 209599) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209600 && (row * 640 + col) <= 209605) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209606 && (row * 640 + col) <= 209611) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209612 && (row * 640 + col) <= 209617) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209618 && (row * 640 + col) <= 209623) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209624 && (row * 640 + col) <= 209629) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209630 && (row * 640 + col) <= 209632) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209633 && (row * 640 + col) <= 209638) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209639 && (row * 640 + col) <= 209641) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209642 && (row * 640 + col) <= 209647) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209648 && (row * 640 + col) <= 209650) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209651 && (row * 640 + col) <= 209656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209657 && (row * 640 + col) <= 209659) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209660 && (row * 640 + col) <= 209665) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209666 && (row * 640 + col) <= 209667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209668 && (row * 640 + col) <= 209680) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209681 && (row * 640 + col) <= 209686) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209687 && (row * 640 + col) <= 209692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209693 && (row * 640 + col) <= 209695) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209696 && (row * 640 + col) <= 209701) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209702 && (row * 640 + col) <= 209707) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209708 && (row * 640 + col) <= 209713) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209714 && (row * 640 + col) <= 209716) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209717 && (row * 640 + col) <= 209722) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209723 && (row * 640 + col) <= 209725) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209726 && (row * 640 + col) <= 209731) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209732 && (row * 640 + col) <= 209737) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209738 && (row * 640 + col) <= 209743) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209744 && (row * 640 + col) <= 209755) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209756 && (row * 640 + col) <= 209761) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209762 && (row * 640 + col) <= 209778) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209779 && (row * 640 + col) <= 209784) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209785 && (row * 640 + col) <= 209807) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209808 && (row * 640 + col) <= 209869) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 209870 && (row * 640 + col) <= 209919) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 209920 && (row * 640 + col) <= 209956) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 209957 && (row * 640 + col) <= 210006) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210007 && (row * 640 + col) <= 210067) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 210068 && (row * 640 + col) <= 210091) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210092 && (row * 640 + col) <= 210109) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210110 && (row * 640 + col) <= 210115) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210116 && (row * 640 + col) <= 210150) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 210151 && (row * 640 + col) <= 210152) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210153 && (row * 640 + col) <= 210155) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210156 && (row * 640 + col) <= 210168) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210169 && (row * 640 + col) <= 210189) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210190 && (row * 640 + col) <= 210197) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210198 && (row * 640 + col) <= 210203) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210204 && (row * 640 + col) <= 210209) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210210 && (row * 640 + col) <= 210215) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210216 && (row * 640 + col) <= 210221) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210222 && (row * 640 + col) <= 210227) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210228 && (row * 640 + col) <= 210239) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210240 && (row * 640 + col) <= 210245) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210246 && (row * 640 + col) <= 210251) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210252 && (row * 640 + col) <= 210257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210258 && (row * 640 + col) <= 210263) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210264 && (row * 640 + col) <= 210269) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210270 && (row * 640 + col) <= 210272) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210273 && (row * 640 + col) <= 210278) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210279 && (row * 640 + col) <= 210281) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210282 && (row * 640 + col) <= 210287) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210288 && (row * 640 + col) <= 210290) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210291 && (row * 640 + col) <= 210296) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210297 && (row * 640 + col) <= 210299) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210300 && (row * 640 + col) <= 210305) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210306 && (row * 640 + col) <= 210307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210308 && (row * 640 + col) <= 210320) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210321 && (row * 640 + col) <= 210326) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210327 && (row * 640 + col) <= 210332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210333 && (row * 640 + col) <= 210335) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210336 && (row * 640 + col) <= 210341) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210342 && (row * 640 + col) <= 210347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210348 && (row * 640 + col) <= 210353) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210354 && (row * 640 + col) <= 210356) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210357 && (row * 640 + col) <= 210362) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210363 && (row * 640 + col) <= 210365) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210366 && (row * 640 + col) <= 210371) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210372 && (row * 640 + col) <= 210377) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210378 && (row * 640 + col) <= 210383) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210384 && (row * 640 + col) <= 210395) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210396 && (row * 640 + col) <= 210401) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210402 && (row * 640 + col) <= 210418) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210419 && (row * 640 + col) <= 210424) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210425 && (row * 640 + col) <= 210447) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210448 && (row * 640 + col) <= 210509) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210510 && (row * 640 + col) <= 210559) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 210560 && (row * 640 + col) <= 210596) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210597 && (row * 640 + col) <= 210645) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210646 && (row * 640 + col) <= 210709) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 210710 && (row * 640 + col) <= 210731) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210732 && (row * 640 + col) <= 210752) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210753 && (row * 640 + col) <= 210758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210759 && (row * 640 + col) <= 210790) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 210791 && (row * 640 + col) <= 210792) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210793 && (row * 640 + col) <= 210795) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210796 && (row * 640 + col) <= 210808) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210809 && (row * 640 + col) <= 210829) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210830 && (row * 640 + col) <= 210837) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210838 && (row * 640 + col) <= 210843) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210844 && (row * 640 + col) <= 210849) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210850 && (row * 640 + col) <= 210855) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210856 && (row * 640 + col) <= 210861) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210862 && (row * 640 + col) <= 210867) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210868 && (row * 640 + col) <= 210879) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210880 && (row * 640 + col) <= 210885) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210886 && (row * 640 + col) <= 210891) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210892 && (row * 640 + col) <= 210897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210898 && (row * 640 + col) <= 210903) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210904 && (row * 640 + col) <= 210909) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210910 && (row * 640 + col) <= 210912) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210913 && (row * 640 + col) <= 210918) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210919 && (row * 640 + col) <= 210921) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210922 && (row * 640 + col) <= 210927) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210928 && (row * 640 + col) <= 210930) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210931 && (row * 640 + col) <= 210936) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210937 && (row * 640 + col) <= 210939) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210940 && (row * 640 + col) <= 210945) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210946 && (row * 640 + col) <= 210947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210948 && (row * 640 + col) <= 210960) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210961 && (row * 640 + col) <= 210966) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210967 && (row * 640 + col) <= 210972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 210973 && (row * 640 + col) <= 210975) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210976 && (row * 640 + col) <= 210981) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210982 && (row * 640 + col) <= 210987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210988 && (row * 640 + col) <= 210993) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210994 && (row * 640 + col) <= 210996) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 210997 && (row * 640 + col) <= 211002) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211003 && (row * 640 + col) <= 211005) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211006 && (row * 640 + col) <= 211011) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211012 && (row * 640 + col) <= 211017) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211018 && (row * 640 + col) <= 211023) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211024 && (row * 640 + col) <= 211035) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211036 && (row * 640 + col) <= 211041) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211042 && (row * 640 + col) <= 211058) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211059 && (row * 640 + col) <= 211064) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211065 && (row * 640 + col) <= 211087) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211088 && (row * 640 + col) <= 211144) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211145 && (row * 640 + col) <= 211199) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 211200 && (row * 640 + col) <= 211236) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211237 && (row * 640 + col) <= 211284) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211285 && (row * 640 + col) <= 211349) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 211350 && (row * 640 + col) <= 211371) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211372 && (row * 640 + col) <= 211394) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211395 && (row * 640 + col) <= 211400) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211401 && (row * 640 + col) <= 211431) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 211432 && (row * 640 + col) <= 211433) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211434 && (row * 640 + col) <= 211435) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211436 && (row * 640 + col) <= 211448) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211449 && (row * 640 + col) <= 211469) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211470 && (row * 640 + col) <= 211477) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211478 && (row * 640 + col) <= 211483) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211484 && (row * 640 + col) <= 211489) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211490 && (row * 640 + col) <= 211495) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211496 && (row * 640 + col) <= 211501) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211502 && (row * 640 + col) <= 211507) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211508 && (row * 640 + col) <= 211519) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211520 && (row * 640 + col) <= 211525) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211526 && (row * 640 + col) <= 211531) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211532 && (row * 640 + col) <= 211537) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211538 && (row * 640 + col) <= 211543) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211544 && (row * 640 + col) <= 211549) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211550 && (row * 640 + col) <= 211552) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211553 && (row * 640 + col) <= 211558) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211559 && (row * 640 + col) <= 211561) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211562 && (row * 640 + col) <= 211567) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211568 && (row * 640 + col) <= 211570) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211571 && (row * 640 + col) <= 211576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211577 && (row * 640 + col) <= 211579) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211580 && (row * 640 + col) <= 211585) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211586 && (row * 640 + col) <= 211587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211588 && (row * 640 + col) <= 211600) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211601 && (row * 640 + col) <= 211606) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211607 && (row * 640 + col) <= 211612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211613 && (row * 640 + col) <= 211615) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211616 && (row * 640 + col) <= 211621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211622 && (row * 640 + col) <= 211627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211628 && (row * 640 + col) <= 211633) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211634 && (row * 640 + col) <= 211636) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211637 && (row * 640 + col) <= 211642) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211643 && (row * 640 + col) <= 211645) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211646 && (row * 640 + col) <= 211651) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211652 && (row * 640 + col) <= 211657) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211658 && (row * 640 + col) <= 211663) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211664 && (row * 640 + col) <= 211675) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211676 && (row * 640 + col) <= 211681) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211682 && (row * 640 + col) <= 211698) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211699 && (row * 640 + col) <= 211704) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211705 && (row * 640 + col) <= 211727) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211728 && (row * 640 + col) <= 211783) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211784 && (row * 640 + col) <= 211817) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 211818 && (row * 640 + col) <= 211826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211827 && (row * 640 + col) <= 211839) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 211840 && (row * 640 + col) <= 211876) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 211877 && (row * 640 + col) <= 211922) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211923 && (row * 640 + col) <= 211989) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 211990 && (row * 640 + col) <= 211992) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 211993 && (row * 640 + col) <= 211994) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 211995 && (row * 640 + col) <= 212011) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212012 && (row * 640 + col) <= 212037) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212038 && (row * 640 + col) <= 212042) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212043 && (row * 640 + col) <= 212071) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 212072 && (row * 640 + col) <= 212073) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212074 && (row * 640 + col) <= 212075) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212076 && (row * 640 + col) <= 212088) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212089 && (row * 640 + col) <= 212109) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212110 && (row * 640 + col) <= 212117) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212118 && (row * 640 + col) <= 212123) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212124 && (row * 640 + col) <= 212129) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212130 && (row * 640 + col) <= 212135) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212136 && (row * 640 + col) <= 212141) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212142 && (row * 640 + col) <= 212147) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212148 && (row * 640 + col) <= 212159) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212160 && (row * 640 + col) <= 212165) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212166 && (row * 640 + col) <= 212171) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212172 && (row * 640 + col) <= 212177) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212178 && (row * 640 + col) <= 212183) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212184 && (row * 640 + col) <= 212189) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212190 && (row * 640 + col) <= 212192) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212193 && (row * 640 + col) <= 212198) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212199 && (row * 640 + col) <= 212201) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212202 && (row * 640 + col) <= 212207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212208 && (row * 640 + col) <= 212210) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212211 && (row * 640 + col) <= 212216) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212217 && (row * 640 + col) <= 212219) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212220 && (row * 640 + col) <= 212225) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212226 && (row * 640 + col) <= 212227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212228 && (row * 640 + col) <= 212240) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212241 && (row * 640 + col) <= 212246) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212247 && (row * 640 + col) <= 212252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212253 && (row * 640 + col) <= 212255) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212256 && (row * 640 + col) <= 212261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212262 && (row * 640 + col) <= 212267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212268 && (row * 640 + col) <= 212273) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212274 && (row * 640 + col) <= 212276) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212277 && (row * 640 + col) <= 212282) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212283 && (row * 640 + col) <= 212285) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212286 && (row * 640 + col) <= 212291) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212292 && (row * 640 + col) <= 212297) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212298 && (row * 640 + col) <= 212303) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212304 && (row * 640 + col) <= 212315) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212316 && (row * 640 + col) <= 212321) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212322 && (row * 640 + col) <= 212338) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212339 && (row * 640 + col) <= 212344) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212345 && (row * 640 + col) <= 212367) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212368 && (row * 640 + col) <= 212423) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212424 && (row * 640 + col) <= 212457) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 212458 && (row * 640 + col) <= 212467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212468 && (row * 640 + col) <= 212479) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 212480 && (row * 640 + col) <= 212517) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212518 && (row * 640 + col) <= 212562) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212563 && (row * 640 + col) <= 212635) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 212636 && (row * 640 + col) <= 212651) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212652 && (row * 640 + col) <= 212677) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212678 && (row * 640 + col) <= 212679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212680 && (row * 640 + col) <= 212684) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212685 && (row * 640 + col) <= 212712) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 212713 && (row * 640 + col) <= 212714) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212715 && (row * 640 + col) <= 212715) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212716 && (row * 640 + col) <= 212728) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212729 && (row * 640 + col) <= 212731) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212732 && (row * 640 + col) <= 212735) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212736 && (row * 640 + col) <= 212736) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 212737 && (row * 640 + col) <= 212749) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212750 && (row * 640 + col) <= 212757) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212758 && (row * 640 + col) <= 212763) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212764 && (row * 640 + col) <= 212769) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212770 && (row * 640 + col) <= 212775) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212776 && (row * 640 + col) <= 212781) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212782 && (row * 640 + col) <= 212787) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212788 && (row * 640 + col) <= 212799) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212800 && (row * 640 + col) <= 212805) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212806 && (row * 640 + col) <= 212811) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212812 && (row * 640 + col) <= 212817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212818 && (row * 640 + col) <= 212823) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212824 && (row * 640 + col) <= 212829) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212830 && (row * 640 + col) <= 212832) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212833 && (row * 640 + col) <= 212838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212839 && (row * 640 + col) <= 212841) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212842 && (row * 640 + col) <= 212847) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212848 && (row * 640 + col) <= 212850) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212851 && (row * 640 + col) <= 212856) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212857 && (row * 640 + col) <= 212859) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212860 && (row * 640 + col) <= 212865) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212866 && (row * 640 + col) <= 212867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212868 && (row * 640 + col) <= 212880) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212881 && (row * 640 + col) <= 212886) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212887 && (row * 640 + col) <= 212892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212893 && (row * 640 + col) <= 212895) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212896 && (row * 640 + col) <= 212901) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212902 && (row * 640 + col) <= 212907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212908 && (row * 640 + col) <= 212913) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212914 && (row * 640 + col) <= 212916) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212917 && (row * 640 + col) <= 212922) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212923 && (row * 640 + col) <= 212925) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212926 && (row * 640 + col) <= 212931) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212932 && (row * 640 + col) <= 212937) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212938 && (row * 640 + col) <= 212943) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212944 && (row * 640 + col) <= 212955) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212956 && (row * 640 + col) <= 212961) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212962 && (row * 640 + col) <= 212978) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 212979 && (row * 640 + col) <= 212984) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 212985 && (row * 640 + col) <= 213007) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213008 && (row * 640 + col) <= 213064) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213065 && (row * 640 + col) <= 213096) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213097 && (row * 640 + col) <= 213107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213108 && (row * 640 + col) <= 213119) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213120 && (row * 640 + col) <= 213165) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213166 && (row * 640 + col) <= 213201) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213202 && (row * 640 + col) <= 213257) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213258 && (row * 640 + col) <= 213271) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213272 && (row * 640 + col) <= 213275) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213276 && (row * 640 + col) <= 213291) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213292 && (row * 640 + col) <= 213317) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213318 && (row * 640 + col) <= 213321) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213322 && (row * 640 + col) <= 213326) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213327 && (row * 640 + col) <= 213352) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 213353 && (row * 640 + col) <= 213354) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213355 && (row * 640 + col) <= 213355) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213356 && (row * 640 + col) <= 213368) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213369 && (row * 640 + col) <= 213371) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213372 && (row * 640 + col) <= 213375) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213376 && (row * 640 + col) <= 213389) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213390 && (row * 640 + col) <= 213397) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213398 && (row * 640 + col) <= 213403) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213404 && (row * 640 + col) <= 213409) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213410 && (row * 640 + col) <= 213415) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213416 && (row * 640 + col) <= 213421) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213422 && (row * 640 + col) <= 213427) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213428 && (row * 640 + col) <= 213430) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213431 && (row * 640 + col) <= 213436) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213437 && (row * 640 + col) <= 213439) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213440 && (row * 640 + col) <= 213445) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213446 && (row * 640 + col) <= 213451) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213452 && (row * 640 + col) <= 213457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213458 && (row * 640 + col) <= 213463) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213464 && (row * 640 + col) <= 213469) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213470 && (row * 640 + col) <= 213472) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213473 && (row * 640 + col) <= 213478) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213479 && (row * 640 + col) <= 213481) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213482 && (row * 640 + col) <= 213487) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213488 && (row * 640 + col) <= 213490) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213491 && (row * 640 + col) <= 213496) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213497 && (row * 640 + col) <= 213499) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213500 && (row * 640 + col) <= 213505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213506 && (row * 640 + col) <= 213507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213508 && (row * 640 + col) <= 213508) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213509 && (row * 640 + col) <= 213514) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213515 && (row * 640 + col) <= 213520) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213521 && (row * 640 + col) <= 213526) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213527 && (row * 640 + col) <= 213532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213533 && (row * 640 + col) <= 213535) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213536 && (row * 640 + col) <= 213541) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213542 && (row * 640 + col) <= 213547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213548 && (row * 640 + col) <= 213553) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213554 && (row * 640 + col) <= 213556) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213557 && (row * 640 + col) <= 213562) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213563 && (row * 640 + col) <= 213565) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213566 && (row * 640 + col) <= 213571) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213572 && (row * 640 + col) <= 213577) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213578 && (row * 640 + col) <= 213583) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213584 && (row * 640 + col) <= 213586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213587 && (row * 640 + col) <= 213592) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213593 && (row * 640 + col) <= 213595) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213596 && (row * 640 + col) <= 213601) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213602 && (row * 640 + col) <= 213618) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213619 && (row * 640 + col) <= 213624) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213625 && (row * 640 + col) <= 213647) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213648 && (row * 640 + col) <= 213704) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213705 && (row * 640 + col) <= 213706) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213707 && (row * 640 + col) <= 213749) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213750 && (row * 640 + col) <= 213750) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213751 && (row * 640 + col) <= 213759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213760 && (row * 640 + col) <= 213805) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213806 && (row * 640 + col) <= 213836) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213837 && (row * 640 + col) <= 213897) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213898 && (row * 640 + col) <= 213911) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213912 && (row * 640 + col) <= 213915) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 213916 && (row * 640 + col) <= 213931) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213932 && (row * 640 + col) <= 213957) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 213958 && (row * 640 + col) <= 213963) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213964 && (row * 640 + col) <= 213968) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213969 && (row * 640 + col) <= 213992) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 213993 && (row * 640 + col) <= 213994) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213995 && (row * 640 + col) <= 213995) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 213996 && (row * 640 + col) <= 214008) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214009 && (row * 640 + col) <= 214011) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214012 && (row * 640 + col) <= 214015) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214016 && (row * 640 + col) <= 214029) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214030 && (row * 640 + col) <= 214037) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214038 && (row * 640 + col) <= 214043) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214044 && (row * 640 + col) <= 214049) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214050 && (row * 640 + col) <= 214055) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214056 && (row * 640 + col) <= 214061) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214062 && (row * 640 + col) <= 214067) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214068 && (row * 640 + col) <= 214070) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214071 && (row * 640 + col) <= 214076) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214077 && (row * 640 + col) <= 214079) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214080 && (row * 640 + col) <= 214085) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214086 && (row * 640 + col) <= 214091) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214092 && (row * 640 + col) <= 214097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214098 && (row * 640 + col) <= 214103) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214104 && (row * 640 + col) <= 214109) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214110 && (row * 640 + col) <= 214112) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214113 && (row * 640 + col) <= 214118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214119 && (row * 640 + col) <= 214121) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214122 && (row * 640 + col) <= 214127) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214128 && (row * 640 + col) <= 214130) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214131 && (row * 640 + col) <= 214136) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214137 && (row * 640 + col) <= 214139) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214140 && (row * 640 + col) <= 214145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214146 && (row * 640 + col) <= 214147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214148 && (row * 640 + col) <= 214148) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214149 && (row * 640 + col) <= 214154) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214155 && (row * 640 + col) <= 214160) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214161 && (row * 640 + col) <= 214166) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214167 && (row * 640 + col) <= 214172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214173 && (row * 640 + col) <= 214175) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214176 && (row * 640 + col) <= 214181) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214182 && (row * 640 + col) <= 214187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214188 && (row * 640 + col) <= 214193) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214194 && (row * 640 + col) <= 214196) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214197 && (row * 640 + col) <= 214202) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214203 && (row * 640 + col) <= 214205) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214206 && (row * 640 + col) <= 214211) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214212 && (row * 640 + col) <= 214217) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214218 && (row * 640 + col) <= 214223) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214224 && (row * 640 + col) <= 214226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214227 && (row * 640 + col) <= 214232) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214233 && (row * 640 + col) <= 214235) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214236 && (row * 640 + col) <= 214241) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214242 && (row * 640 + col) <= 214258) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214259 && (row * 640 + col) <= 214264) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214265 && (row * 640 + col) <= 214287) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214288 && (row * 640 + col) <= 214399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214400 && (row * 640 + col) <= 214445) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214446 && (row * 640 + col) <= 214475) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214476 && (row * 640 + col) <= 214537) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 214538 && (row * 640 + col) <= 214605) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214606 && (row * 640 + col) <= 214610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214611 && (row * 640 + col) <= 214632) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 214633 && (row * 640 + col) <= 214634) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214635 && (row * 640 + col) <= 214648) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214649 && (row * 640 + col) <= 214651) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214652 && (row * 640 + col) <= 214655) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214656 && (row * 640 + col) <= 214669) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214670 && (row * 640 + col) <= 214677) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214678 && (row * 640 + col) <= 214683) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214684 && (row * 640 + col) <= 214689) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214690 && (row * 640 + col) <= 214695) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214696 && (row * 640 + col) <= 214701) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214702 && (row * 640 + col) <= 214707) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214708 && (row * 640 + col) <= 214710) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214711 && (row * 640 + col) <= 214716) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214717 && (row * 640 + col) <= 214719) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214720 && (row * 640 + col) <= 214725) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214726 && (row * 640 + col) <= 214731) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214732 && (row * 640 + col) <= 214737) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214738 && (row * 640 + col) <= 214743) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214744 && (row * 640 + col) <= 214749) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214750 && (row * 640 + col) <= 214752) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214753 && (row * 640 + col) <= 214758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214759 && (row * 640 + col) <= 214761) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214762 && (row * 640 + col) <= 214767) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214768 && (row * 640 + col) <= 214770) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214771 && (row * 640 + col) <= 214776) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214777 && (row * 640 + col) <= 214779) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214780 && (row * 640 + col) <= 214785) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214786 && (row * 640 + col) <= 214787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214788 && (row * 640 + col) <= 214788) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214789 && (row * 640 + col) <= 214794) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214795 && (row * 640 + col) <= 214800) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214801 && (row * 640 + col) <= 214806) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214807 && (row * 640 + col) <= 214812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214813 && (row * 640 + col) <= 214815) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214816 && (row * 640 + col) <= 214821) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214822 && (row * 640 + col) <= 214827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214828 && (row * 640 + col) <= 214833) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214834 && (row * 640 + col) <= 214836) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214837 && (row * 640 + col) <= 214842) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214843 && (row * 640 + col) <= 214845) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214846 && (row * 640 + col) <= 214851) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214852 && (row * 640 + col) <= 214857) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214858 && (row * 640 + col) <= 214863) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214864 && (row * 640 + col) <= 214866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214867 && (row * 640 + col) <= 214872) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214873 && (row * 640 + col) <= 214875) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214876 && (row * 640 + col) <= 214881) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214882 && (row * 640 + col) <= 214898) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214899 && (row * 640 + col) <= 214904) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 214905 && (row * 640 + col) <= 214927) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 214928 && (row * 640 + col) <= 215039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215040 && (row * 640 + col) <= 215085) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215086 && (row * 640 + col) <= 215115) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215116 && (row * 640 + col) <= 215177) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 215178 && (row * 640 + col) <= 215247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215248 && (row * 640 + col) <= 215251) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215252 && (row * 640 + col) <= 215272) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 215273 && (row * 640 + col) <= 215274) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215275 && (row * 640 + col) <= 215288) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215289 && (row * 640 + col) <= 215309) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215310 && (row * 640 + col) <= 215314) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215315 && (row * 640 + col) <= 215326) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215327 && (row * 640 + col) <= 215329) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215330 && (row * 640 + col) <= 215335) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215336 && (row * 640 + col) <= 215341) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215342 && (row * 640 + col) <= 215347) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215348 && (row * 640 + col) <= 215350) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215351 && (row * 640 + col) <= 215365) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215366 && (row * 640 + col) <= 215371) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215372 && (row * 640 + col) <= 215377) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215378 && (row * 640 + col) <= 215383) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215384 && (row * 640 + col) <= 215389) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215390 && (row * 640 + col) <= 215392) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215393 && (row * 640 + col) <= 215398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215399 && (row * 640 + col) <= 215401) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215402 && (row * 640 + col) <= 215416) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215417 && (row * 640 + col) <= 215419) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215420 && (row * 640 + col) <= 215434) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215435 && (row * 640 + col) <= 215440) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215441 && (row * 640 + col) <= 215446) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215447 && (row * 640 + col) <= 215452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215453 && (row * 640 + col) <= 215464) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215465 && (row * 640 + col) <= 215467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215468 && (row * 640 + col) <= 215482) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215483 && (row * 640 + col) <= 215485) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215486 && (row * 640 + col) <= 215491) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215492 && (row * 640 + col) <= 215497) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215498 && (row * 640 + col) <= 215503) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215504 && (row * 640 + col) <= 215506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215507 && (row * 640 + col) <= 215521) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215522 && (row * 640 + col) <= 215538) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215539 && (row * 640 + col) <= 215544) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215545 && (row * 640 + col) <= 215567) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215568 && (row * 640 + col) <= 215679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215680 && (row * 640 + col) <= 215725) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215726 && (row * 640 + col) <= 215754) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215755 && (row * 640 + col) <= 215817) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 215818 && (row * 640 + col) <= 215889) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215890 && (row * 640 + col) <= 215892) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215893 && (row * 640 + col) <= 215912) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 215913 && (row * 640 + col) <= 215914) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215915 && (row * 640 + col) <= 215928) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215929 && (row * 640 + col) <= 215949) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215950 && (row * 640 + col) <= 215954) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215955 && (row * 640 + col) <= 215966) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215967 && (row * 640 + col) <= 215969) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215970 && (row * 640 + col) <= 215975) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215976 && (row * 640 + col) <= 215981) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 215982 && (row * 640 + col) <= 215987) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215988 && (row * 640 + col) <= 215990) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 215991 && (row * 640 + col) <= 216005) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216006 && (row * 640 + col) <= 216011) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216012 && (row * 640 + col) <= 216017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216018 && (row * 640 + col) <= 216023) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216024 && (row * 640 + col) <= 216029) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216030 && (row * 640 + col) <= 216032) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216033 && (row * 640 + col) <= 216038) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216039 && (row * 640 + col) <= 216041) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216042 && (row * 640 + col) <= 216056) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216057 && (row * 640 + col) <= 216059) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216060 && (row * 640 + col) <= 216074) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216075 && (row * 640 + col) <= 216080) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216081 && (row * 640 + col) <= 216086) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216087 && (row * 640 + col) <= 216092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216093 && (row * 640 + col) <= 216104) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216105 && (row * 640 + col) <= 216107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216108 && (row * 640 + col) <= 216122) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216123 && (row * 640 + col) <= 216125) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216126 && (row * 640 + col) <= 216131) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216132 && (row * 640 + col) <= 216137) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216138 && (row * 640 + col) <= 216143) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216144 && (row * 640 + col) <= 216146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216147 && (row * 640 + col) <= 216161) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216162 && (row * 640 + col) <= 216178) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216179 && (row * 640 + col) <= 216184) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216185 && (row * 640 + col) <= 216207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216208 && (row * 640 + col) <= 216319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216320 && (row * 640 + col) <= 216365) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216366 && (row * 640 + col) <= 216390) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216391 && (row * 640 + col) <= 216457) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 216458 && (row * 640 + col) <= 216530) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216531 && (row * 640 + col) <= 216534) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216535 && (row * 640 + col) <= 216551) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 216552 && (row * 640 + col) <= 216554) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216555 && (row * 640 + col) <= 216555) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216556 && (row * 640 + col) <= 216568) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216569 && (row * 640 + col) <= 216589) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216590 && (row * 640 + col) <= 216594) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216595 && (row * 640 + col) <= 216606) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216607 && (row * 640 + col) <= 216609) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216610 && (row * 640 + col) <= 216615) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216616 && (row * 640 + col) <= 216621) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216622 && (row * 640 + col) <= 216627) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216628 && (row * 640 + col) <= 216630) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216631 && (row * 640 + col) <= 216645) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216646 && (row * 640 + col) <= 216651) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216652 && (row * 640 + col) <= 216657) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216658 && (row * 640 + col) <= 216663) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216664 && (row * 640 + col) <= 216669) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216670 && (row * 640 + col) <= 216672) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216673 && (row * 640 + col) <= 216678) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216679 && (row * 640 + col) <= 216681) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216682 && (row * 640 + col) <= 216696) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216697 && (row * 640 + col) <= 216699) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216700 && (row * 640 + col) <= 216714) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216715 && (row * 640 + col) <= 216720) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216721 && (row * 640 + col) <= 216726) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216727 && (row * 640 + col) <= 216732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216733 && (row * 640 + col) <= 216744) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216745 && (row * 640 + col) <= 216747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216748 && (row * 640 + col) <= 216762) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216763 && (row * 640 + col) <= 216765) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216766 && (row * 640 + col) <= 216771) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216772 && (row * 640 + col) <= 216777) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216778 && (row * 640 + col) <= 216783) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216784 && (row * 640 + col) <= 216786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216787 && (row * 640 + col) <= 216801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216802 && (row * 640 + col) <= 216818) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216819 && (row * 640 + col) <= 216824) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216825 && (row * 640 + col) <= 216847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 216848 && (row * 640 + col) <= 216959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 216960 && (row * 640 + col) <= 217005) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217006 && (row * 640 + col) <= 217030) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217031 && (row * 640 + col) <= 217097) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 217098 && (row * 640 + col) <= 217171) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217172 && (row * 640 + col) <= 217176) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217177 && (row * 640 + col) <= 217191) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 217192 && (row * 640 + col) <= 217193) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217194 && (row * 640 + col) <= 217195) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217196 && (row * 640 + col) <= 217208) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217209 && (row * 640 + col) <= 217229) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217230 && (row * 640 + col) <= 217251) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217252 && (row * 640 + col) <= 217266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217267 && (row * 640 + col) <= 217295) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217296 && (row * 640 + col) <= 217306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217307 && (row * 640 + col) <= 217332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217333 && (row * 640 + col) <= 217347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217348 && (row * 640 + col) <= 217372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217373 && (row * 640 + col) <= 217441) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217442 && (row * 640 + col) <= 217458) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217459 && (row * 640 + col) <= 217464) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217465 && (row * 640 + col) <= 217487) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217488 && (row * 640 + col) <= 217599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217600 && (row * 640 + col) <= 217645) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217646 && (row * 640 + col) <= 217665) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217666 && (row * 640 + col) <= 217737) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 217738 && (row * 640 + col) <= 217813) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217814 && (row * 640 + col) <= 217818) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217819 && (row * 640 + col) <= 217830) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 217831 && (row * 640 + col) <= 217833) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217834 && (row * 640 + col) <= 217835) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217836 && (row * 640 + col) <= 217848) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217849 && (row * 640 + col) <= 217869) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217870 && (row * 640 + col) <= 217891) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217892 && (row * 640 + col) <= 217906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217907 && (row * 640 + col) <= 217935) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217936 && (row * 640 + col) <= 217946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217947 && (row * 640 + col) <= 217972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 217973 && (row * 640 + col) <= 217987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 217988 && (row * 640 + col) <= 218012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218013 && (row * 640 + col) <= 218081) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218082 && (row * 640 + col) <= 218098) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218099 && (row * 640 + col) <= 218104) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218105 && (row * 640 + col) <= 218127) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218128 && (row * 640 + col) <= 218239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218240 && (row * 640 + col) <= 218285) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218286 && (row * 640 + col) <= 218304) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218305 && (row * 640 + col) <= 218377) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 218378 && (row * 640 + col) <= 218455) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218456 && (row * 640 + col) <= 218460) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218461 && (row * 640 + col) <= 218469) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 218470 && (row * 640 + col) <= 218472) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218473 && (row * 640 + col) <= 218475) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218476 && (row * 640 + col) <= 218488) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218489 && (row * 640 + col) <= 218509) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218510 && (row * 640 + col) <= 218531) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218532 && (row * 640 + col) <= 218546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218547 && (row * 640 + col) <= 218577) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218578 && (row * 640 + col) <= 218583) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218584 && (row * 640 + col) <= 218612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218613 && (row * 640 + col) <= 218627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218628 && (row * 640 + col) <= 218661) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218662 && (row * 640 + col) <= 218721) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218722 && (row * 640 + col) <= 218738) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218739 && (row * 640 + col) <= 218744) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218745 && (row * 640 + col) <= 218767) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218768 && (row * 640 + col) <= 218879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218880 && (row * 640 + col) <= 218925) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 218926 && (row * 640 + col) <= 218943) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 218944 && (row * 640 + col) <= 219017) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 219018 && (row * 640 + col) <= 219097) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219098 && (row * 640 + col) <= 219102) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219103 && (row * 640 + col) <= 219107) color_data <= 12'b011000101111; else
        if ((row * 640 + col) >= 219108 && (row * 640 + col) <= 219111) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219112 && (row * 640 + col) <= 219115) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219116 && (row * 640 + col) <= 219128) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219129 && (row * 640 + col) <= 219149) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219150 && (row * 640 + col) <= 219171) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219172 && (row * 640 + col) <= 219186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219187 && (row * 640 + col) <= 219217) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219218 && (row * 640 + col) <= 219223) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219224 && (row * 640 + col) <= 219252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219253 && (row * 640 + col) <= 219267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219268 && (row * 640 + col) <= 219301) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219302 && (row * 640 + col) <= 219361) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219362 && (row * 640 + col) <= 219378) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219379 && (row * 640 + col) <= 219384) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219385 && (row * 640 + col) <= 219407) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219408 && (row * 640 + col) <= 219519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219520 && (row * 640 + col) <= 219565) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219566 && (row * 640 + col) <= 219581) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219582 && (row * 640 + col) <= 219657) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 219658 && (row * 640 + col) <= 219739) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219740 && (row * 640 + col) <= 219750) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219751 && (row * 640 + col) <= 219755) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219756 && (row * 640 + col) <= 219768) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219769 && (row * 640 + col) <= 219789) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219790 && (row * 640 + col) <= 219811) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219812 && (row * 640 + col) <= 219826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219827 && (row * 640 + col) <= 219857) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219858 && (row * 640 + col) <= 219863) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219864 && (row * 640 + col) <= 219892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219893 && (row * 640 + col) <= 219907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 219908 && (row * 640 + col) <= 219941) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 219942 && (row * 640 + col) <= 220001) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220002 && (row * 640 + col) <= 220018) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220019 && (row * 640 + col) <= 220024) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220025 && (row * 640 + col) <= 220047) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220048 && (row * 640 + col) <= 220159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220160 && (row * 640 + col) <= 220205) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220206 && (row * 640 + col) <= 220221) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220222 && (row * 640 + col) <= 220297) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 220298 && (row * 640 + col) <= 220381) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220382 && (row * 640 + col) <= 220388) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220389 && (row * 640 + col) <= 220395) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220396 && (row * 640 + col) <= 220408) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220409 && (row * 640 + col) <= 220429) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220430 && (row * 640 + col) <= 220451) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220452 && (row * 640 + col) <= 220466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220467 && (row * 640 + col) <= 220497) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220498 && (row * 640 + col) <= 220503) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220504 && (row * 640 + col) <= 220532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220533 && (row * 640 + col) <= 220547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220548 && (row * 640 + col) <= 220581) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220582 && (row * 640 + col) <= 220641) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220642 && (row * 640 + col) <= 220658) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220659 && (row * 640 + col) <= 220664) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220665 && (row * 640 + col) <= 220687) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220688 && (row * 640 + col) <= 220799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220800 && (row * 640 + col) <= 220845) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 220846 && (row * 640 + col) <= 220860) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 220861 && (row * 640 + col) <= 220937) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 220938 && (row * 640 + col) <= 221028) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221029 && (row * 640 + col) <= 221035) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221036 && (row * 640 + col) <= 221048) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221049 && (row * 640 + col) <= 221069) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221070 && (row * 640 + col) <= 221091) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221092 && (row * 640 + col) <= 221106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221107 && (row * 640 + col) <= 221137) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221138 && (row * 640 + col) <= 221143) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221144 && (row * 640 + col) <= 221172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221173 && (row * 640 + col) <= 221187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221188 && (row * 640 + col) <= 221221) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221222 && (row * 640 + col) <= 221281) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221282 && (row * 640 + col) <= 221298) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221299 && (row * 640 + col) <= 221304) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221305 && (row * 640 + col) <= 221327) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221328 && (row * 640 + col) <= 221439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221440 && (row * 640 + col) <= 221485) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221486 && (row * 640 + col) <= 221496) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221497 && (row * 640 + col) <= 221576) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 221577 && (row * 640 + col) <= 221577) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221578 && (row * 640 + col) <= 221668) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221669 && (row * 640 + col) <= 221674) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221675 && (row * 640 + col) <= 221688) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221689 && (row * 640 + col) <= 221709) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221710 && (row * 640 + col) <= 221732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221733 && (row * 640 + col) <= 221746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221747 && (row * 640 + col) <= 221777) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221778 && (row * 640 + col) <= 221783) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221784 && (row * 640 + col) <= 221812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221813 && (row * 640 + col) <= 221827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221828 && (row * 640 + col) <= 221861) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221862 && (row * 640 + col) <= 221921) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221922 && (row * 640 + col) <= 221938) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221939 && (row * 640 + col) <= 221944) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 221945 && (row * 640 + col) <= 221967) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 221968 && (row * 640 + col) <= 222079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222080 && (row * 640 + col) <= 222125) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222126 && (row * 640 + col) <= 222135) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222136 && (row * 640 + col) <= 222215) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 222216 && (row * 640 + col) <= 222217) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222218 && (row * 640 + col) <= 222328) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222329 && (row * 640 + col) <= 222349) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222350 && (row * 640 + col) <= 222380) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222381 && (row * 640 + col) <= 222386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222387 && (row * 640 + col) <= 222417) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222418 && (row * 640 + col) <= 222423) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222424 && (row * 640 + col) <= 222452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222453 && (row * 640 + col) <= 222467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222468 && (row * 640 + col) <= 222501) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222502 && (row * 640 + col) <= 222561) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222562 && (row * 640 + col) <= 222607) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222608 && (row * 640 + col) <= 222719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222720 && (row * 640 + col) <= 222765) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222766 && (row * 640 + col) <= 222775) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222776 && (row * 640 + col) <= 222787) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 222788 && (row * 640 + col) <= 222790) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222791 && (row * 640 + col) <= 222809) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 222810 && (row * 640 + col) <= 222821) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222822 && (row * 640 + col) <= 222841) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 222842 && (row * 640 + col) <= 222857) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222858 && (row * 640 + col) <= 222968) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 222969 && (row * 640 + col) <= 222989) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 222990 && (row * 640 + col) <= 223020) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223021 && (row * 640 + col) <= 223026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223027 && (row * 640 + col) <= 223057) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223058 && (row * 640 + col) <= 223063) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223064 && (row * 640 + col) <= 223092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223093 && (row * 640 + col) <= 223107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223108 && (row * 640 + col) <= 223141) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223142 && (row * 640 + col) <= 223201) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223202 && (row * 640 + col) <= 223247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223248 && (row * 640 + col) <= 223359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223360 && (row * 640 + col) <= 223405) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223406 && (row * 640 + col) <= 223415) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223416 && (row * 640 + col) <= 223426) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 223427 && (row * 640 + col) <= 223430) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223431 && (row * 640 + col) <= 223449) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 223450 && (row * 640 + col) <= 223461) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223462 && (row * 640 + col) <= 223481) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 223482 && (row * 640 + col) <= 223497) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223498 && (row * 640 + col) <= 223608) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223609 && (row * 640 + col) <= 223629) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223630 && (row * 640 + col) <= 223660) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223661 && (row * 640 + col) <= 223666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223667 && (row * 640 + col) <= 223697) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223698 && (row * 640 + col) <= 223703) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223704 && (row * 640 + col) <= 223732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223733 && (row * 640 + col) <= 223747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223748 && (row * 640 + col) <= 223781) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223782 && (row * 640 + col) <= 223841) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 223842 && (row * 640 + col) <= 223887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 223888 && (row * 640 + col) <= 223999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224000 && (row * 640 + col) <= 224045) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224046 && (row * 640 + col) <= 224058) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224059 && (row * 640 + col) <= 224059) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 224060 && (row * 640 + col) <= 224103) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224104 && (row * 640 + col) <= 224104) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 224105 && (row * 640 + col) <= 224112) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224113 && (row * 640 + col) <= 224113) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 224114 && (row * 640 + col) <= 224137) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224138 && (row * 640 + col) <= 224248) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224249 && (row * 640 + col) <= 224269) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224270 && (row * 640 + col) <= 224300) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224301 && (row * 640 + col) <= 224306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224307 && (row * 640 + col) <= 224337) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224338 && (row * 640 + col) <= 224343) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224344 && (row * 640 + col) <= 224372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224373 && (row * 640 + col) <= 224387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224388 && (row * 640 + col) <= 224421) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224422 && (row * 640 + col) <= 224481) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224482 && (row * 640 + col) <= 224527) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224528 && (row * 640 + col) <= 224639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224640 && (row * 640 + col) <= 224685) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224686 && (row * 640 + col) <= 224777) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224778 && (row * 640 + col) <= 224888) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224889 && (row * 640 + col) <= 224909) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224910 && (row * 640 + col) <= 224940) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224941 && (row * 640 + col) <= 224946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224947 && (row * 640 + col) <= 224977) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 224978 && (row * 640 + col) <= 224983) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 224984 && (row * 640 + col) <= 225012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225013 && (row * 640 + col) <= 225027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225028 && (row * 640 + col) <= 225061) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225062 && (row * 640 + col) <= 225121) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225122 && (row * 640 + col) <= 225167) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225168 && (row * 640 + col) <= 225279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225280 && (row * 640 + col) <= 225325) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225326 && (row * 640 + col) <= 225354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225355 && (row * 640 + col) <= 225358) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225359 && (row * 640 + col) <= 225364) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225365 && (row * 640 + col) <= 225367) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225368 && (row * 640 + col) <= 225381) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225382 && (row * 640 + col) <= 225382) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225383 && (row * 640 + col) <= 225383) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225384 && (row * 640 + col) <= 225384) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225385 && (row * 640 + col) <= 225417) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225418 && (row * 640 + col) <= 225528) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225529 && (row * 640 + col) <= 225549) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225550 && (row * 640 + col) <= 225580) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225581 && (row * 640 + col) <= 225586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225587 && (row * 640 + col) <= 225617) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225618 && (row * 640 + col) <= 225623) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225624 && (row * 640 + col) <= 225652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225653 && (row * 640 + col) <= 225667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225668 && (row * 640 + col) <= 225701) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225702 && (row * 640 + col) <= 225708) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225709 && (row * 640 + col) <= 225728) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225729 && (row * 640 + col) <= 225729) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225730 && (row * 640 + col) <= 225732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225733 && (row * 640 + col) <= 225743) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225744 && (row * 640 + col) <= 225745) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225746 && (row * 640 + col) <= 225747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225748 && (row * 640 + col) <= 225749) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225750 && (row * 640 + col) <= 225750) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225751 && (row * 640 + col) <= 225807) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225808 && (row * 640 + col) <= 225919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225920 && (row * 640 + col) <= 225965) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 225966 && (row * 640 + col) <= 225994) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 225995 && (row * 640 + col) <= 226025) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226026 && (row * 640 + col) <= 226057) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226058 && (row * 640 + col) <= 226168) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226169 && (row * 640 + col) <= 226189) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226190 && (row * 640 + col) <= 226220) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226221 && (row * 640 + col) <= 226226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226227 && (row * 640 + col) <= 226257) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226258 && (row * 640 + col) <= 226263) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226264 && (row * 640 + col) <= 226292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226293 && (row * 640 + col) <= 226307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226308 && (row * 640 + col) <= 226341) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226342 && (row * 640 + col) <= 226347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226348 && (row * 640 + col) <= 226372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226373 && (row * 640 + col) <= 226381) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226382 && (row * 640 + col) <= 226447) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226448 && (row * 640 + col) <= 226559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226560 && (row * 640 + col) <= 226605) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226606 && (row * 640 + col) <= 226634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226635 && (row * 640 + col) <= 226665) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226666 && (row * 640 + col) <= 226697) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226698 && (row * 640 + col) <= 226808) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226809 && (row * 640 + col) <= 226829) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226830 && (row * 640 + col) <= 226860) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226861 && (row * 640 + col) <= 226866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226867 && (row * 640 + col) <= 226897) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226898 && (row * 640 + col) <= 226903) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226904 && (row * 640 + col) <= 226932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226933 && (row * 640 + col) <= 226947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226948 && (row * 640 + col) <= 226981) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 226982 && (row * 640 + col) <= 226987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 226988 && (row * 640 + col) <= 227012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227013 && (row * 640 + col) <= 227021) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227022 && (row * 640 + col) <= 227087) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227088 && (row * 640 + col) <= 227199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227200 && (row * 640 + col) <= 227245) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227246 && (row * 640 + col) <= 227274) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227275 && (row * 640 + col) <= 227305) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227306 && (row * 640 + col) <= 227337) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227338 && (row * 640 + col) <= 227449) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227450 && (row * 640 + col) <= 227450) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227451 && (row * 640 + col) <= 227451) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227452 && (row * 640 + col) <= 227469) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227470 && (row * 640 + col) <= 227500) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227501 && (row * 640 + col) <= 227506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227507 && (row * 640 + col) <= 227537) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227538 && (row * 640 + col) <= 227541) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227542 && (row * 640 + col) <= 227542) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227543 && (row * 640 + col) <= 227543) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227544 && (row * 640 + col) <= 227572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227573 && (row * 640 + col) <= 227587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227588 && (row * 640 + col) <= 227621) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227622 && (row * 640 + col) <= 227627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227628 && (row * 640 + col) <= 227652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227653 && (row * 640 + col) <= 227661) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227662 && (row * 640 + col) <= 227727) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227728 && (row * 640 + col) <= 227839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227840 && (row * 640 + col) <= 227885) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227886 && (row * 640 + col) <= 227914) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227915 && (row * 640 + col) <= 227945) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 227946 && (row * 640 + col) <= 227977) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 227978 && (row * 640 + col) <= 228091) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228092 && (row * 640 + col) <= 228109) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228110 && (row * 640 + col) <= 228140) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228141 && (row * 640 + col) <= 228146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228147 && (row * 640 + col) <= 228177) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228178 && (row * 640 + col) <= 228181) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228182 && (row * 640 + col) <= 228212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228213 && (row * 640 + col) <= 228227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228228 && (row * 640 + col) <= 228261) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228262 && (row * 640 + col) <= 228267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228268 && (row * 640 + col) <= 228292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228293 && (row * 640 + col) <= 228301) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228302 && (row * 640 + col) <= 228367) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228368 && (row * 640 + col) <= 228479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228480 && (row * 640 + col) <= 228525) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228526 && (row * 640 + col) <= 228554) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228555 && (row * 640 + col) <= 228585) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228586 && (row * 640 + col) <= 228617) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228618 && (row * 640 + col) <= 228731) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228732 && (row * 640 + col) <= 228749) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228750 && (row * 640 + col) <= 228780) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228781 && (row * 640 + col) <= 228786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228787 && (row * 640 + col) <= 228817) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228818 && (row * 640 + col) <= 228821) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228822 && (row * 640 + col) <= 228852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228853 && (row * 640 + col) <= 228867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228868 && (row * 640 + col) <= 228901) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228902 && (row * 640 + col) <= 228907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228908 && (row * 640 + col) <= 228932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 228933 && (row * 640 + col) <= 228941) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 228942 && (row * 640 + col) <= 229007) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229008 && (row * 640 + col) <= 229119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229120 && (row * 640 + col) <= 229165) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229166 && (row * 640 + col) <= 229194) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229195 && (row * 640 + col) <= 229225) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229226 && (row * 640 + col) <= 229257) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229258 && (row * 640 + col) <= 229371) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229372 && (row * 640 + col) <= 229389) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229390 && (row * 640 + col) <= 229420) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229421 && (row * 640 + col) <= 229426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229427 && (row * 640 + col) <= 229457) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229458 && (row * 640 + col) <= 229461) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229462 && (row * 640 + col) <= 229541) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229542 && (row * 640 + col) <= 229547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229548 && (row * 640 + col) <= 229572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229573 && (row * 640 + col) <= 229581) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229582 && (row * 640 + col) <= 229647) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229648 && (row * 640 + col) <= 229759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229760 && (row * 640 + col) <= 229805) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229806 && (row * 640 + col) <= 229834) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229835 && (row * 640 + col) <= 229865) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 229866 && (row * 640 + col) <= 229897) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 229898 && (row * 640 + col) <= 230011) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230012 && (row * 640 + col) <= 230029) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230030 && (row * 640 + col) <= 230060) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230061 && (row * 640 + col) <= 230066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230067 && (row * 640 + col) <= 230097) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230098 && (row * 640 + col) <= 230101) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230102 && (row * 640 + col) <= 230181) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230182 && (row * 640 + col) <= 230187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230188 && (row * 640 + col) <= 230212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230213 && (row * 640 + col) <= 230221) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230222 && (row * 640 + col) <= 230287) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230288 && (row * 640 + col) <= 230399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230400 && (row * 640 + col) <= 230445) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230446 && (row * 640 + col) <= 230474) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230475 && (row * 640 + col) <= 230505) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230506 && (row * 640 + col) <= 230537) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230538 && (row * 640 + col) <= 230651) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230652 && (row * 640 + col) <= 230669) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230670 && (row * 640 + col) <= 230700) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230701 && (row * 640 + col) <= 230706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230707 && (row * 640 + col) <= 230737) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230738 && (row * 640 + col) <= 230741) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230742 && (row * 640 + col) <= 230821) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230822 && (row * 640 + col) <= 230827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230828 && (row * 640 + col) <= 230852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230853 && (row * 640 + col) <= 230861) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 230862 && (row * 640 + col) <= 230927) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 230928 && (row * 640 + col) <= 231039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231040 && (row * 640 + col) <= 231085) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231086 && (row * 640 + col) <= 231111) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231112 && (row * 640 + col) <= 231148) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231149 && (row * 640 + col) <= 231177) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231178 && (row * 640 + col) <= 231291) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231292 && (row * 640 + col) <= 231309) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231310 && (row * 640 + col) <= 231340) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231341 && (row * 640 + col) <= 231346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231347 && (row * 640 + col) <= 231461) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231462 && (row * 640 + col) <= 231467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231468 && (row * 640 + col) <= 231492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231493 && (row * 640 + col) <= 231501) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231502 && (row * 640 + col) <= 231567) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231568 && (row * 640 + col) <= 231679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231680 && (row * 640 + col) <= 231725) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231726 && (row * 640 + col) <= 231751) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231752 && (row * 640 + col) <= 231788) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231789 && (row * 640 + col) <= 231817) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231818 && (row * 640 + col) <= 231931) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231932 && (row * 640 + col) <= 231949) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231950 && (row * 640 + col) <= 231980) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 231981 && (row * 640 + col) <= 231986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 231987 && (row * 640 + col) <= 232101) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232102 && (row * 640 + col) <= 232107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232108 && (row * 640 + col) <= 232132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232133 && (row * 640 + col) <= 232141) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232142 && (row * 640 + col) <= 232207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232208 && (row * 640 + col) <= 232319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232320 && (row * 640 + col) <= 232365) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232366 && (row * 640 + col) <= 232391) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232392 && (row * 640 + col) <= 232428) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232429 && (row * 640 + col) <= 232457) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232458 && (row * 640 + col) <= 232571) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232572 && (row * 640 + col) <= 232589) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232590 && (row * 640 + col) <= 232620) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232621 && (row * 640 + col) <= 232626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232627 && (row * 640 + col) <= 232741) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232742 && (row * 640 + col) <= 232747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232748 && (row * 640 + col) <= 232772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232773 && (row * 640 + col) <= 232781) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232782 && (row * 640 + col) <= 232847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 232848 && (row * 640 + col) <= 232959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 232960 && (row * 640 + col) <= 233005) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233006 && (row * 640 + col) <= 233031) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233032 && (row * 640 + col) <= 233068) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233069 && (row * 640 + col) <= 233097) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233098 && (row * 640 + col) <= 233211) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233212 && (row * 640 + col) <= 233220) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233221 && (row * 640 + col) <= 233226) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233227 && (row * 640 + col) <= 233229) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233230 && (row * 640 + col) <= 233263) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233264 && (row * 640 + col) <= 233266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233267 && (row * 640 + col) <= 233381) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233382 && (row * 640 + col) <= 233387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233388 && (row * 640 + col) <= 233412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233413 && (row * 640 + col) <= 233421) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233422 && (row * 640 + col) <= 233487) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233488 && (row * 640 + col) <= 233599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233600 && (row * 640 + col) <= 233645) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233646 && (row * 640 + col) <= 233671) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233672 && (row * 640 + col) <= 233708) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233709 && (row * 640 + col) <= 233737) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233738 && (row * 640 + col) <= 233851) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233852 && (row * 640 + col) <= 233860) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233861 && (row * 640 + col) <= 233866) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233867 && (row * 640 + col) <= 233869) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233870 && (row * 640 + col) <= 233903) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 233904 && (row * 640 + col) <= 233906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 233907 && (row * 640 + col) <= 234021) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234022 && (row * 640 + col) <= 234027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234028 && (row * 640 + col) <= 234052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234053 && (row * 640 + col) <= 234061) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234062 && (row * 640 + col) <= 234127) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234128 && (row * 640 + col) <= 234239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234240 && (row * 640 + col) <= 234285) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234286 && (row * 640 + col) <= 234311) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234312 && (row * 640 + col) <= 234348) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234349 && (row * 640 + col) <= 234377) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234378 && (row * 640 + col) <= 234491) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234492 && (row * 640 + col) <= 234500) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234501 && (row * 640 + col) <= 234506) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234507 && (row * 640 + col) <= 234509) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234510 && (row * 640 + col) <= 234543) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234544 && (row * 640 + col) <= 234546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234547 && (row * 640 + col) <= 234661) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234662 && (row * 640 + col) <= 234667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234668 && (row * 640 + col) <= 234692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234693 && (row * 640 + col) <= 234701) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234702 && (row * 640 + col) <= 234767) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234768 && (row * 640 + col) <= 234879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234880 && (row * 640 + col) <= 234925) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234926 && (row * 640 + col) <= 234951) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 234952 && (row * 640 + col) <= 234988) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 234989 && (row * 640 + col) <= 235017) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235018 && (row * 640 + col) <= 235131) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235132 && (row * 640 + col) <= 235138) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235139 && (row * 640 + col) <= 235183) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235184 && (row * 640 + col) <= 235186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235187 && (row * 640 + col) <= 235301) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235302 && (row * 640 + col) <= 235307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235308 && (row * 640 + col) <= 235332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235333 && (row * 640 + col) <= 235341) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235342 && (row * 640 + col) <= 235407) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235408 && (row * 640 + col) <= 235519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235520 && (row * 640 + col) <= 235565) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235566 && (row * 640 + col) <= 235591) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235592 && (row * 640 + col) <= 235628) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235629 && (row * 640 + col) <= 235657) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235658 && (row * 640 + col) <= 235771) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235772 && (row * 640 + col) <= 235777) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235778 && (row * 640 + col) <= 235823) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235824 && (row * 640 + col) <= 235826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235827 && (row * 640 + col) <= 235941) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235942 && (row * 640 + col) <= 235947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235948 && (row * 640 + col) <= 235972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 235973 && (row * 640 + col) <= 235981) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 235982 && (row * 640 + col) <= 236047) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236048 && (row * 640 + col) <= 236159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236160 && (row * 640 + col) <= 236205) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236206 && (row * 640 + col) <= 236231) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236232 && (row * 640 + col) <= 236268) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236269 && (row * 640 + col) <= 236297) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236298 && (row * 640 + col) <= 236411) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236412 && (row * 640 + col) <= 236417) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236418 && (row * 640 + col) <= 236463) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236464 && (row * 640 + col) <= 236466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236467 && (row * 640 + col) <= 236581) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236582 && (row * 640 + col) <= 236587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236588 && (row * 640 + col) <= 236612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236613 && (row * 640 + col) <= 236621) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236622 && (row * 640 + col) <= 236687) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236688 && (row * 640 + col) <= 236738) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236739 && (row * 640 + col) <= 236748) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 236749 && (row * 640 + col) <= 236799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236800 && (row * 640 + col) <= 236845) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236846 && (row * 640 + col) <= 236871) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236872 && (row * 640 + col) <= 236908) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236909 && (row * 640 + col) <= 236920) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236921 && (row * 640 + col) <= 236928) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 236929 && (row * 640 + col) <= 236937) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 236938 && (row * 640 + col) <= 237103) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237104 && (row * 640 + col) <= 237106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237107 && (row * 640 + col) <= 237221) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237222 && (row * 640 + col) <= 237227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237228 && (row * 640 + col) <= 237327) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237328 && (row * 640 + col) <= 237378) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237379 && (row * 640 + col) <= 237389) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 237390 && (row * 640 + col) <= 237439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237440 && (row * 640 + col) <= 237485) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237486 && (row * 640 + col) <= 237511) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237512 && (row * 640 + col) <= 237548) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237549 && (row * 640 + col) <= 237560) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237561 && (row * 640 + col) <= 237568) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237569 && (row * 640 + col) <= 237577) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237578 && (row * 640 + col) <= 237743) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237744 && (row * 640 + col) <= 237746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237747 && (row * 640 + col) <= 237861) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237862 && (row * 640 + col) <= 237867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 237868 && (row * 640 + col) <= 237967) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 237968 && (row * 640 + col) <= 238017) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238018 && (row * 640 + col) <= 238029) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 238030 && (row * 640 + col) <= 238033) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238034 && (row * 640 + col) <= 238036) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 238037 && (row * 640 + col) <= 238079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238080 && (row * 640 + col) <= 238125) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238126 && (row * 640 + col) <= 238151) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238152 && (row * 640 + col) <= 238188) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238189 && (row * 640 + col) <= 238199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238200 && (row * 640 + col) <= 238208) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238209 && (row * 640 + col) <= 238217) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238218 && (row * 640 + col) <= 238383) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238384 && (row * 640 + col) <= 238386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238387 && (row * 640 + col) <= 238501) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238502 && (row * 640 + col) <= 238507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238508 && (row * 640 + col) <= 238607) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238608 && (row * 640 + col) <= 238655) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238656 && (row * 640 + col) <= 238677) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 238678 && (row * 640 + col) <= 238719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238720 && (row * 640 + col) <= 238765) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238766 && (row * 640 + col) <= 238788) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238789 && (row * 640 + col) <= 238828) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 238829 && (row * 640 + col) <= 238831) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 238832 && (row * 640 + col) <= 239141) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239142 && (row * 640 + col) <= 239147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239148 && (row * 640 + col) <= 239247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239248 && (row * 640 + col) <= 239262) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239263 && (row * 640 + col) <= 239267) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239268 && (row * 640 + col) <= 239295) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239296 && (row * 640 + col) <= 239317) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 239318 && (row * 640 + col) <= 239359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239360 && (row * 640 + col) <= 239405) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239406 && (row * 640 + col) <= 239428) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239429 && (row * 640 + col) <= 239468) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239469 && (row * 640 + col) <= 239471) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239472 && (row * 640 + col) <= 239781) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239782 && (row * 640 + col) <= 239787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239788 && (row * 640 + col) <= 239887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239888 && (row * 640 + col) <= 239902) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239903 && (row * 640 + col) <= 239907) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 239908 && (row * 640 + col) <= 239934) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 239935 && (row * 640 + col) <= 239958) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 239959 && (row * 640 + col) <= 239999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240000 && (row * 640 + col) <= 240045) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240046 && (row * 640 + col) <= 240068) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240069 && (row * 640 + col) <= 240108) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240109 && (row * 640 + col) <= 240111) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240112 && (row * 640 + col) <= 240195) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240196 && (row * 640 + col) <= 240212) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240213 && (row * 640 + col) <= 240421) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240422 && (row * 640 + col) <= 240427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240428 && (row * 640 + col) <= 240527) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240528 && (row * 640 + col) <= 240541) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240542 && (row * 640 + col) <= 240548) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240549 && (row * 640 + col) <= 240572) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240573 && (row * 640 + col) <= 240600) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 240601 && (row * 640 + col) <= 240639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240640 && (row * 640 + col) <= 240685) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240686 && (row * 640 + col) <= 240708) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240709 && (row * 640 + col) <= 240748) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240749 && (row * 640 + col) <= 240751) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 240752 && (row * 640 + col) <= 240828) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 240829 && (row * 640 + col) <= 240857) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240858 && (row * 640 + col) <= 241061) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241062 && (row * 640 + col) <= 241067) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241068 && (row * 640 + col) <= 241196) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241197 && (row * 640 + col) <= 241212) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241213 && (row * 640 + col) <= 241240) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 241241 && (row * 640 + col) <= 241279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241280 && (row * 640 + col) <= 241325) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241326 && (row * 640 + col) <= 241348) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241349 && (row * 640 + col) <= 241388) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241389 && (row * 640 + col) <= 241391) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241392 && (row * 640 + col) <= 241462) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241463 && (row * 640 + col) <= 241476) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241477 && (row * 640 + col) <= 241491) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241492 && (row * 640 + col) <= 241501) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241502 && (row * 640 + col) <= 241701) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241702 && (row * 640 + col) <= 241707) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241708 && (row * 640 + col) <= 241836) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241837 && (row * 640 + col) <= 241839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241840 && (row * 640 + col) <= 241880) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 241881 && (row * 640 + col) <= 241919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241920 && (row * 640 + col) <= 241965) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 241966 && (row * 640 + col) <= 241988) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 241989 && (row * 640 + col) <= 242028) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242029 && (row * 640 + col) <= 242031) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 242032 && (row * 640 + col) <= 242099) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242100 && (row * 640 + col) <= 242109) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242110 && (row * 640 + col) <= 242136) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242137 && (row * 640 + col) <= 242143) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242144 && (row * 640 + col) <= 242341) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242342 && (row * 640 + col) <= 242347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 242348 && (row * 640 + col) <= 242476) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242477 && (row * 640 + col) <= 242478) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 242479 && (row * 640 + col) <= 242520) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 242521 && (row * 640 + col) <= 242559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 242560 && (row * 640 + col) <= 242605) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242606 && (row * 640 + col) <= 242628) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 242629 && (row * 640 + col) <= 242668) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242669 && (row * 640 + col) <= 242671) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 242672 && (row * 640 + col) <= 242736) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242737 && (row * 640 + col) <= 242743) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242744 && (row * 640 + col) <= 242780) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242781 && (row * 640 + col) <= 242786) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242787 && (row * 640 + col) <= 242981) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 242982 && (row * 640 + col) <= 242987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 242988 && (row * 640 + col) <= 243116) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243117 && (row * 640 + col) <= 243118) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243119 && (row * 640 + col) <= 243160) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 243161 && (row * 640 + col) <= 243199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243200 && (row * 640 + col) <= 243245) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243246 && (row * 640 + col) <= 243268) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243269 && (row * 640 + col) <= 243308) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243309 && (row * 640 + col) <= 243311) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243312 && (row * 640 + col) <= 243373) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243374 && (row * 640 + col) <= 243380) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243381 && (row * 640 + col) <= 243422) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243423 && (row * 640 + col) <= 243428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243429 && (row * 640 + col) <= 243621) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243622 && (row * 640 + col) <= 243627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243628 && (row * 640 + col) <= 243756) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243757 && (row * 640 + col) <= 243804) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 243805 && (row * 640 + col) <= 243839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243840 && (row * 640 + col) <= 243890) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243891 && (row * 640 + col) <= 243899) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243900 && (row * 640 + col) <= 243948) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 243949 && (row * 640 + col) <= 243951) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 243952 && (row * 640 + col) <= 244011) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 244012 && (row * 640 + col) <= 244017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244018 && (row * 640 + col) <= 244065) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244066 && (row * 640 + col) <= 244069) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244070 && (row * 640 + col) <= 244261) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 244262 && (row * 640 + col) <= 244267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 244268 && (row * 640 + col) <= 244396) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 244397 && (row * 640 + col) <= 244445) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 244446 && (row * 640 + col) <= 244479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 244480 && (row * 640 + col) <= 244530) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 244531 && (row * 640 + col) <= 244539) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 244540 && (row * 640 + col) <= 244588) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 244589 && (row * 640 + col) <= 244591) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 244592 && (row * 640 + col) <= 244648) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 244649 && (row * 640 + col) <= 244654) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244655 && (row * 640 + col) <= 244707) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244708 && (row * 640 + col) <= 244711) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244712 && (row * 640 + col) <= 244901) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 244902 && (row * 640 + col) <= 244907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 244908 && (row * 640 + col) <= 245036) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245037 && (row * 640 + col) <= 245086) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 245087 && (row * 640 + col) <= 245119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 245120 && (row * 640 + col) <= 245170) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245171 && (row * 640 + col) <= 245179) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 245180 && (row * 640 + col) <= 245228) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245229 && (row * 640 + col) <= 245231) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 245232 && (row * 640 + col) <= 245287) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245288 && (row * 640 + col) <= 245292) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245293 && (row * 640 + col) <= 245349) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245350 && (row * 640 + col) <= 245352) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245353 && (row * 640 + col) <= 245541) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245542 && (row * 640 + col) <= 245547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 245548 && (row * 640 + col) <= 245676) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245677 && (row * 640 + col) <= 245730) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 245731 && (row * 640 + col) <= 245759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 245760 && (row * 640 + col) <= 245810) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245811 && (row * 640 + col) <= 245819) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 245820 && (row * 640 + col) <= 245868) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245869 && (row * 640 + col) <= 245871) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 245872 && (row * 640 + col) <= 245925) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 245926 && (row * 640 + col) <= 245929) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245930 && (row * 640 + col) <= 245990) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245991 && (row * 640 + col) <= 245993) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245994 && (row * 640 + col) <= 246316) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 246317 && (row * 640 + col) <= 246371) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 246372 && (row * 640 + col) <= 246399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 246400 && (row * 640 + col) <= 246450) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 246451 && (row * 640 + col) <= 246459) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 246460 && (row * 640 + col) <= 246508) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 246509 && (row * 640 + col) <= 246511) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 246512 && (row * 640 + col) <= 246563) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 246564 && (row * 640 + col) <= 246568) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246569 && (row * 640 + col) <= 246631) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246632 && (row * 640 + col) <= 246634) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246635 && (row * 640 + col) <= 246956) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 246957 && (row * 640 + col) <= 247011) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 247012 && (row * 640 + col) <= 247039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 247040 && (row * 640 + col) <= 247090) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247091 && (row * 640 + col) <= 247099) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 247100 && (row * 640 + col) <= 247148) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247149 && (row * 640 + col) <= 247151) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 247152 && (row * 640 + col) <= 247202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247203 && (row * 640 + col) <= 247206) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247207 && (row * 640 + col) <= 247272) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247273 && (row * 640 + col) <= 247274) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247275 && (row * 640 + col) <= 247312) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247313 && (row * 640 + col) <= 247324) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247325 && (row * 640 + col) <= 247327) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247328 && (row * 640 + col) <= 247342) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247343 && (row * 640 + col) <= 247345) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247346 && (row * 640 + col) <= 247360) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247361 && (row * 640 + col) <= 247363) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247364 && (row * 640 + col) <= 247375) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247376 && (row * 640 + col) <= 247384) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247385 && (row * 640 + col) <= 247399) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247400 && (row * 640 + col) <= 247402) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247403 && (row * 640 + col) <= 247417) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247418 && (row * 640 + col) <= 247420) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247421 && (row * 640 + col) <= 247426) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247427 && (row * 640 + col) <= 247432) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247433 && (row * 640 + col) <= 247438) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247439 && (row * 640 + col) <= 247441) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247442 && (row * 640 + col) <= 247453) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247454 && (row * 640 + col) <= 247456) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247457 && (row * 640 + col) <= 247471) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247472 && (row * 640 + col) <= 247474) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247475 && (row * 640 + col) <= 247489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247490 && (row * 640 + col) <= 247492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247493 && (row * 640 + col) <= 247498) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247499 && (row * 640 + col) <= 247510) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247511 && (row * 640 + col) <= 247516) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247517 && (row * 640 + col) <= 247528) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247529 && (row * 640 + col) <= 247543) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247544 && (row * 640 + col) <= 247546) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247547 && (row * 640 + col) <= 247561) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247562 && (row * 640 + col) <= 247596) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247597 && (row * 640 + col) <= 247651) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 247652 && (row * 640 + col) <= 247679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 247680 && (row * 640 + col) <= 247730) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247731 && (row * 640 + col) <= 247739) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 247740 && (row * 640 + col) <= 247788) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247789 && (row * 640 + col) <= 247791) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 247792 && (row * 640 + col) <= 247840) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247841 && (row * 640 + col) <= 247844) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247845 && (row * 640 + col) <= 247865) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247866 && (row * 640 + col) <= 247871) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247872 && (row * 640 + col) <= 247874) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247875 && (row * 640 + col) <= 247880) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247881 && (row * 640 + col) <= 247913) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247914 && (row * 640 + col) <= 247915) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247916 && (row * 640 + col) <= 247952) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247953 && (row * 640 + col) <= 247964) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247965 && (row * 640 + col) <= 247967) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247968 && (row * 640 + col) <= 247982) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247983 && (row * 640 + col) <= 247985) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 247986 && (row * 640 + col) <= 248000) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248001 && (row * 640 + col) <= 248003) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248004 && (row * 640 + col) <= 248015) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248016 && (row * 640 + col) <= 248024) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248025 && (row * 640 + col) <= 248039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248040 && (row * 640 + col) <= 248042) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248043 && (row * 640 + col) <= 248057) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248058 && (row * 640 + col) <= 248060) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248061 && (row * 640 + col) <= 248066) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248067 && (row * 640 + col) <= 248072) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248073 && (row * 640 + col) <= 248078) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248079 && (row * 640 + col) <= 248081) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248082 && (row * 640 + col) <= 248093) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248094 && (row * 640 + col) <= 248096) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248097 && (row * 640 + col) <= 248111) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248112 && (row * 640 + col) <= 248114) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248115 && (row * 640 + col) <= 248129) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248130 && (row * 640 + col) <= 248132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248133 && (row * 640 + col) <= 248138) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248139 && (row * 640 + col) <= 248150) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248151 && (row * 640 + col) <= 248156) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248157 && (row * 640 + col) <= 248168) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248169 && (row * 640 + col) <= 248183) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248184 && (row * 640 + col) <= 248186) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248187 && (row * 640 + col) <= 248201) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248202 && (row * 640 + col) <= 248236) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248237 && (row * 640 + col) <= 248237) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 248238 && (row * 640 + col) <= 248290) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 248291 && (row * 640 + col) <= 248319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 248320 && (row * 640 + col) <= 248370) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248371 && (row * 640 + col) <= 248379) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 248380 && (row * 640 + col) <= 248428) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248429 && (row * 640 + col) <= 248431) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 248432 && (row * 640 + col) <= 248479) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248480 && (row * 640 + col) <= 248483) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248484 && (row * 640 + col) <= 248505) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248506 && (row * 640 + col) <= 248511) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248512 && (row * 640 + col) <= 248514) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248515 && (row * 640 + col) <= 248520) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248521 && (row * 640 + col) <= 248553) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248554 && (row * 640 + col) <= 248556) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248557 && (row * 640 + col) <= 248592) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248593 && (row * 640 + col) <= 248604) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248605 && (row * 640 + col) <= 248607) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248608 && (row * 640 + col) <= 248622) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248623 && (row * 640 + col) <= 248625) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248626 && (row * 640 + col) <= 248640) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248641 && (row * 640 + col) <= 248643) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248644 && (row * 640 + col) <= 248655) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248656 && (row * 640 + col) <= 248664) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248665 && (row * 640 + col) <= 248679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248680 && (row * 640 + col) <= 248682) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248683 && (row * 640 + col) <= 248697) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248698 && (row * 640 + col) <= 248700) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248701 && (row * 640 + col) <= 248706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248707 && (row * 640 + col) <= 248712) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248713 && (row * 640 + col) <= 248718) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248719 && (row * 640 + col) <= 248721) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248722 && (row * 640 + col) <= 248733) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248734 && (row * 640 + col) <= 248736) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248737 && (row * 640 + col) <= 248751) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248752 && (row * 640 + col) <= 248754) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248755 && (row * 640 + col) <= 248769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248770 && (row * 640 + col) <= 248772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248773 && (row * 640 + col) <= 248778) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248779 && (row * 640 + col) <= 248790) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248791 && (row * 640 + col) <= 248796) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248797 && (row * 640 + col) <= 248808) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248809 && (row * 640 + col) <= 248823) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248824 && (row * 640 + col) <= 248826) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248827 && (row * 640 + col) <= 248841) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248842 && (row * 640 + col) <= 248876) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 248877 && (row * 640 + col) <= 248959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 248960 && (row * 640 + col) <= 249010) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249011 && (row * 640 + col) <= 249019) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 249020 && (row * 640 + col) <= 249068) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249069 && (row * 640 + col) <= 249071) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 249072 && (row * 640 + col) <= 249118) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249119 && (row * 640 + col) <= 249121) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249122 && (row * 640 + col) <= 249145) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 249146 && (row * 640 + col) <= 249151) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249152 && (row * 640 + col) <= 249154) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 249155 && (row * 640 + col) <= 249160) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249161 && (row * 640 + col) <= 249194) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 249195 && (row * 640 + col) <= 249196) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249197 && (row * 640 + col) <= 249209) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249210 && (row * 640 + col) <= 249213) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249214 && (row * 640 + col) <= 249235) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249236 && (row * 640 + col) <= 249241) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249242 && (row * 640 + col) <= 249247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249248 && (row * 640 + col) <= 249253) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249254 && (row * 640 + col) <= 249256) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249257 && (row * 640 + col) <= 249262) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249263 && (row * 640 + col) <= 249265) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249266 && (row * 640 + col) <= 249271) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249272 && (row * 640 + col) <= 249274) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249275 && (row * 640 + col) <= 249280) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249281 && (row * 640 + col) <= 249286) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249287 && (row * 640 + col) <= 249292) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249293 && (row * 640 + col) <= 249304) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249305 && (row * 640 + col) <= 249310) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249311 && (row * 640 + col) <= 249313) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249314 && (row * 640 + col) <= 249319) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249320 && (row * 640 + col) <= 249322) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249323 && (row * 640 + col) <= 249328) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249329 && (row * 640 + col) <= 249331) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249332 && (row * 640 + col) <= 249337) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249338 && (row * 640 + col) <= 249340) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249341 && (row * 640 + col) <= 249349) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249350 && (row * 640 + col) <= 249352) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249353 && (row * 640 + col) <= 249358) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249359 && (row * 640 + col) <= 249364) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249365 && (row * 640 + col) <= 249370) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249371 && (row * 640 + col) <= 249376) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249377 && (row * 640 + col) <= 249382) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249383 && (row * 640 + col) <= 249385) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249386 && (row * 640 + col) <= 249391) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249392 && (row * 640 + col) <= 249394) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249395 && (row * 640 + col) <= 249400) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249401 && (row * 640 + col) <= 249403) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249404 && (row * 640 + col) <= 249409) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249410 && (row * 640 + col) <= 249412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249413 && (row * 640 + col) <= 249418) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249419 && (row * 640 + col) <= 249430) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249431 && (row * 640 + col) <= 249436) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249437 && (row * 640 + col) <= 249448) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249449 && (row * 640 + col) <= 249454) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249455 && (row * 640 + col) <= 249457) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249458 && (row * 640 + col) <= 249463) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249464 && (row * 640 + col) <= 249466) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249467 && (row * 640 + col) <= 249472) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249473 && (row * 640 + col) <= 249475) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249476 && (row * 640 + col) <= 249481) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249482 && (row * 640 + col) <= 249516) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249517 && (row * 640 + col) <= 249599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 249600 && (row * 640 + col) <= 249650) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249651 && (row * 640 + col) <= 249659) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 249660 && (row * 640 + col) <= 249757) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249758 && (row * 640 + col) <= 249760) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249761 && (row * 640 + col) <= 249785) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 249786 && (row * 640 + col) <= 249791) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249792 && (row * 640 + col) <= 249794) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 249795 && (row * 640 + col) <= 249800) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249801 && (row * 640 + col) <= 249834) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 249835 && (row * 640 + col) <= 249837) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249838 && (row * 640 + col) <= 249849) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249850 && (row * 640 + col) <= 249853) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249854 && (row * 640 + col) <= 249875) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249876 && (row * 640 + col) <= 249881) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249882 && (row * 640 + col) <= 249887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249888 && (row * 640 + col) <= 249893) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249894 && (row * 640 + col) <= 249896) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249897 && (row * 640 + col) <= 249902) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249903 && (row * 640 + col) <= 249905) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249906 && (row * 640 + col) <= 249911) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249912 && (row * 640 + col) <= 249914) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249915 && (row * 640 + col) <= 249920) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249921 && (row * 640 + col) <= 249926) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249927 && (row * 640 + col) <= 249932) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249933 && (row * 640 + col) <= 249944) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249945 && (row * 640 + col) <= 249950) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249951 && (row * 640 + col) <= 249953) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249954 && (row * 640 + col) <= 249959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249960 && (row * 640 + col) <= 249962) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249963 && (row * 640 + col) <= 249968) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249969 && (row * 640 + col) <= 249971) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249972 && (row * 640 + col) <= 249977) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249978 && (row * 640 + col) <= 249980) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249981 && (row * 640 + col) <= 249989) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249990 && (row * 640 + col) <= 249992) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 249993 && (row * 640 + col) <= 249998) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249999 && (row * 640 + col) <= 250004) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250005 && (row * 640 + col) <= 250010) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250011 && (row * 640 + col) <= 250016) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250017 && (row * 640 + col) <= 250022) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250023 && (row * 640 + col) <= 250025) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250026 && (row * 640 + col) <= 250031) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250032 && (row * 640 + col) <= 250034) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250035 && (row * 640 + col) <= 250040) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250041 && (row * 640 + col) <= 250043) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250044 && (row * 640 + col) <= 250049) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250050 && (row * 640 + col) <= 250052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250053 && (row * 640 + col) <= 250058) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250059 && (row * 640 + col) <= 250070) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250071 && (row * 640 + col) <= 250076) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250077 && (row * 640 + col) <= 250088) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250089 && (row * 640 + col) <= 250094) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250095 && (row * 640 + col) <= 250097) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250098 && (row * 640 + col) <= 250103) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250104 && (row * 640 + col) <= 250106) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250107 && (row * 640 + col) <= 250112) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250113 && (row * 640 + col) <= 250115) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250116 && (row * 640 + col) <= 250121) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250122 && (row * 640 + col) <= 250156) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250157 && (row * 640 + col) <= 250239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 250240 && (row * 640 + col) <= 250290) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250291 && (row * 640 + col) <= 250299) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 250300 && (row * 640 + col) <= 250396) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250397 && (row * 640 + col) <= 250399) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250400 && (row * 640 + col) <= 250425) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 250426 && (row * 640 + col) <= 250431) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 250432 && (row * 640 + col) <= 250434) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 250435 && (row * 640 + col) <= 250440) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 250441 && (row * 640 + col) <= 250475) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 250476 && (row * 640 + col) <= 250477) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250478 && (row * 640 + col) <= 250489) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250490 && (row * 640 + col) <= 250493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250494 && (row * 640 + col) <= 250515) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250516 && (row * 640 + col) <= 250521) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250522 && (row * 640 + col) <= 250527) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250528 && (row * 640 + col) <= 250533) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250534 && (row * 640 + col) <= 250536) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250537 && (row * 640 + col) <= 250542) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250543 && (row * 640 + col) <= 250545) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250546 && (row * 640 + col) <= 250551) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250552 && (row * 640 + col) <= 250554) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250555 && (row * 640 + col) <= 250560) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250561 && (row * 640 + col) <= 250566) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250567 && (row * 640 + col) <= 250572) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250573 && (row * 640 + col) <= 250584) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250585 && (row * 640 + col) <= 250590) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250591 && (row * 640 + col) <= 250593) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250594 && (row * 640 + col) <= 250599) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250600 && (row * 640 + col) <= 250602) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250603 && (row * 640 + col) <= 250608) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250609 && (row * 640 + col) <= 250611) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250612 && (row * 640 + col) <= 250617) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250618 && (row * 640 + col) <= 250620) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250621 && (row * 640 + col) <= 250629) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250630 && (row * 640 + col) <= 250632) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250633 && (row * 640 + col) <= 250638) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250639 && (row * 640 + col) <= 250644) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250645 && (row * 640 + col) <= 250650) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250651 && (row * 640 + col) <= 250656) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250657 && (row * 640 + col) <= 250662) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250663 && (row * 640 + col) <= 250665) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250666 && (row * 640 + col) <= 250671) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250672 && (row * 640 + col) <= 250674) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250675 && (row * 640 + col) <= 250680) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250681 && (row * 640 + col) <= 250683) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250684 && (row * 640 + col) <= 250689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250690 && (row * 640 + col) <= 250692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250693 && (row * 640 + col) <= 250698) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250699 && (row * 640 + col) <= 250710) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250711 && (row * 640 + col) <= 250716) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250717 && (row * 640 + col) <= 250728) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250729 && (row * 640 + col) <= 250734) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250735 && (row * 640 + col) <= 250737) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250738 && (row * 640 + col) <= 250743) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250744 && (row * 640 + col) <= 250746) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250747 && (row * 640 + col) <= 250752) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250753 && (row * 640 + col) <= 250755) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250756 && (row * 640 + col) <= 250761) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250762 && (row * 640 + col) <= 250796) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250797 && (row * 640 + col) <= 250879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 250880 && (row * 640 + col) <= 250931) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 250932 && (row * 640 + col) <= 250939) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 250940 && (row * 640 + col) <= 251035) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251036 && (row * 640 + col) <= 251038) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251039 && (row * 640 + col) <= 251065) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 251066 && (row * 640 + col) <= 251071) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251072 && (row * 640 + col) <= 251074) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 251075 && (row * 640 + col) <= 251080) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251081 && (row * 640 + col) <= 251116) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 251117 && (row * 640 + col) <= 251118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251119 && (row * 640 + col) <= 251129) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251130 && (row * 640 + col) <= 251133) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251134 && (row * 640 + col) <= 251155) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251156 && (row * 640 + col) <= 251161) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251162 && (row * 640 + col) <= 251167) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251168 && (row * 640 + col) <= 251173) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251174 && (row * 640 + col) <= 251185) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251186 && (row * 640 + col) <= 251191) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251192 && (row * 640 + col) <= 251206) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251207 && (row * 640 + col) <= 251212) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251213 && (row * 640 + col) <= 251224) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251225 && (row * 640 + col) <= 251230) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251231 && (row * 640 + col) <= 251242) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251243 && (row * 640 + col) <= 251248) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251249 && (row * 640 + col) <= 251251) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251252 && (row * 640 + col) <= 251257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251258 && (row * 640 + col) <= 251260) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251261 && (row * 640 + col) <= 251278) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251279 && (row * 640 + col) <= 251284) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251285 && (row * 640 + col) <= 251290) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251291 && (row * 640 + col) <= 251296) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251297 && (row * 640 + col) <= 251302) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251303 && (row * 640 + col) <= 251305) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251306 && (row * 640 + col) <= 251311) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251312 && (row * 640 + col) <= 251314) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251315 && (row * 640 + col) <= 251320) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251321 && (row * 640 + col) <= 251323) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251324 && (row * 640 + col) <= 251329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251330 && (row * 640 + col) <= 251332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251333 && (row * 640 + col) <= 251338) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251339 && (row * 640 + col) <= 251350) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251351 && (row * 640 + col) <= 251356) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251357 && (row * 640 + col) <= 251368) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251369 && (row * 640 + col) <= 251374) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251375 && (row * 640 + col) <= 251386) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251387 && (row * 640 + col) <= 251392) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251393 && (row * 640 + col) <= 251395) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251396 && (row * 640 + col) <= 251401) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251402 && (row * 640 + col) <= 251436) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251437 && (row * 640 + col) <= 251519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 251520 && (row * 640 + col) <= 251674) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251675 && (row * 640 + col) <= 251677) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251678 && (row * 640 + col) <= 251705) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 251706 && (row * 640 + col) <= 251711) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251712 && (row * 640 + col) <= 251714) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 251715 && (row * 640 + col) <= 251720) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251721 && (row * 640 + col) <= 251756) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 251757 && (row * 640 + col) <= 251758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251759 && (row * 640 + col) <= 251795) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251796 && (row * 640 + col) <= 251801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251802 && (row * 640 + col) <= 251807) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251808 && (row * 640 + col) <= 251813) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251814 && (row * 640 + col) <= 251825) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251826 && (row * 640 + col) <= 251831) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251832 && (row * 640 + col) <= 251846) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251847 && (row * 640 + col) <= 251852) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251853 && (row * 640 + col) <= 251864) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251865 && (row * 640 + col) <= 251870) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251871 && (row * 640 + col) <= 251882) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251883 && (row * 640 + col) <= 251888) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251889 && (row * 640 + col) <= 251891) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251892 && (row * 640 + col) <= 251897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251898 && (row * 640 + col) <= 251900) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251901 && (row * 640 + col) <= 251918) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251919 && (row * 640 + col) <= 251924) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251925 && (row * 640 + col) <= 251930) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251931 && (row * 640 + col) <= 251936) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251937 && (row * 640 + col) <= 251942) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251943 && (row * 640 + col) <= 251945) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251946 && (row * 640 + col) <= 251951) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251952 && (row * 640 + col) <= 251954) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251955 && (row * 640 + col) <= 251960) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251961 && (row * 640 + col) <= 251963) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251964 && (row * 640 + col) <= 251969) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251970 && (row * 640 + col) <= 251972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251973 && (row * 640 + col) <= 251978) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251979 && (row * 640 + col) <= 251990) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 251991 && (row * 640 + col) <= 251996) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251997 && (row * 640 + col) <= 252008) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252009 && (row * 640 + col) <= 252014) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252015 && (row * 640 + col) <= 252026) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252027 && (row * 640 + col) <= 252032) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252033 && (row * 640 + col) <= 252035) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252036 && (row * 640 + col) <= 252041) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252042 && (row * 640 + col) <= 252076) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252077 && (row * 640 + col) <= 252125) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 252126 && (row * 640 + col) <= 252127) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252128 && (row * 640 + col) <= 252159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 252160 && (row * 640 + col) <= 252313) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252314 && (row * 640 + col) <= 252316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252317 && (row * 640 + col) <= 252345) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 252346 && (row * 640 + col) <= 252351) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 252352 && (row * 640 + col) <= 252354) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 252355 && (row * 640 + col) <= 252360) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 252361 && (row * 640 + col) <= 252396) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 252397 && (row * 640 + col) <= 252398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252399 && (row * 640 + col) <= 252435) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252436 && (row * 640 + col) <= 252441) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252442 && (row * 640 + col) <= 252447) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252448 && (row * 640 + col) <= 252453) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252454 && (row * 640 + col) <= 252465) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252466 && (row * 640 + col) <= 252471) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252472 && (row * 640 + col) <= 252486) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252487 && (row * 640 + col) <= 252492) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252493 && (row * 640 + col) <= 252504) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252505 && (row * 640 + col) <= 252510) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252511 && (row * 640 + col) <= 252522) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252523 && (row * 640 + col) <= 252528) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252529 && (row * 640 + col) <= 252531) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252532 && (row * 640 + col) <= 252537) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252538 && (row * 640 + col) <= 252540) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252541 && (row * 640 + col) <= 252558) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252559 && (row * 640 + col) <= 252564) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252565 && (row * 640 + col) <= 252570) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252571 && (row * 640 + col) <= 252576) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252577 && (row * 640 + col) <= 252582) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252583 && (row * 640 + col) <= 252585) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252586 && (row * 640 + col) <= 252591) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252592 && (row * 640 + col) <= 252594) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252595 && (row * 640 + col) <= 252600) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252601 && (row * 640 + col) <= 252603) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252604 && (row * 640 + col) <= 252609) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252610 && (row * 640 + col) <= 252612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252613 && (row * 640 + col) <= 252618) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252619 && (row * 640 + col) <= 252630) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252631 && (row * 640 + col) <= 252636) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252637 && (row * 640 + col) <= 252648) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252649 && (row * 640 + col) <= 252654) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252655 && (row * 640 + col) <= 252666) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252667 && (row * 640 + col) <= 252672) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252673 && (row * 640 + col) <= 252675) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252676 && (row * 640 + col) <= 252681) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252682 && (row * 640 + col) <= 252716) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252717 && (row * 640 + col) <= 252765) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 252766 && (row * 640 + col) <= 252767) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252768 && (row * 640 + col) <= 252799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 252800 && (row * 640 + col) <= 252953) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 252954 && (row * 640 + col) <= 252955) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252956 && (row * 640 + col) <= 252985) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 252986 && (row * 640 + col) <= 252991) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 252992 && (row * 640 + col) <= 252994) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 252995 && (row * 640 + col) <= 253000) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 253001 && (row * 640 + col) <= 253037) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 253038 && (row * 640 + col) <= 253039) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253040 && (row * 640 + col) <= 253075) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253076 && (row * 640 + col) <= 253081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253082 && (row * 640 + col) <= 253087) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253088 && (row * 640 + col) <= 253099) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253100 && (row * 640 + col) <= 253108) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253109 && (row * 640 + col) <= 253117) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253118 && (row * 640 + col) <= 253126) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253127 && (row * 640 + col) <= 253132) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253133 && (row * 640 + col) <= 253144) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253145 && (row * 640 + col) <= 253150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253151 && (row * 640 + col) <= 253162) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253163 && (row * 640 + col) <= 253168) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253169 && (row * 640 + col) <= 253171) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253172 && (row * 640 + col) <= 253177) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253178 && (row * 640 + col) <= 253180) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253181 && (row * 640 + col) <= 253186) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253187 && (row * 640 + col) <= 253189) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253190 && (row * 640 + col) <= 253198) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253199 && (row * 640 + col) <= 253204) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253205 && (row * 640 + col) <= 253210) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253211 && (row * 640 + col) <= 253216) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253217 && (row * 640 + col) <= 253228) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253229 && (row * 640 + col) <= 253234) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253235 && (row * 640 + col) <= 253240) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253241 && (row * 640 + col) <= 253243) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253244 && (row * 640 + col) <= 253249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253250 && (row * 640 + col) <= 253252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253253 && (row * 640 + col) <= 253258) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253259 && (row * 640 + col) <= 253270) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253271 && (row * 640 + col) <= 253276) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253277 && (row * 640 + col) <= 253288) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253289 && (row * 640 + col) <= 253300) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253301 && (row * 640 + col) <= 253306) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253307 && (row * 640 + col) <= 253318) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253319 && (row * 640 + col) <= 253356) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253357 && (row * 640 + col) <= 253404) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 253405 && (row * 640 + col) <= 253408) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253409 && (row * 640 + col) <= 253439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 253440 && (row * 640 + col) <= 253592) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253593 && (row * 640 + col) <= 253595) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253596 && (row * 640 + col) <= 253628) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 253629 && (row * 640 + col) <= 253640) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 253641 && (row * 640 + col) <= 253677) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 253678 && (row * 640 + col) <= 253679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253680 && (row * 640 + col) <= 253715) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253716 && (row * 640 + col) <= 253721) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253722 && (row * 640 + col) <= 253727) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253728 && (row * 640 + col) <= 253739) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253740 && (row * 640 + col) <= 253748) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253749 && (row * 640 + col) <= 253757) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253758 && (row * 640 + col) <= 253766) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253767 && (row * 640 + col) <= 253772) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253773 && (row * 640 + col) <= 253784) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253785 && (row * 640 + col) <= 253790) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253791 && (row * 640 + col) <= 253802) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253803 && (row * 640 + col) <= 253808) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253809 && (row * 640 + col) <= 253811) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253812 && (row * 640 + col) <= 253817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253818 && (row * 640 + col) <= 253820) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253821 && (row * 640 + col) <= 253826) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253827 && (row * 640 + col) <= 253829) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253830 && (row * 640 + col) <= 253838) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253839 && (row * 640 + col) <= 253844) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253845 && (row * 640 + col) <= 253850) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253851 && (row * 640 + col) <= 253856) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253857 && (row * 640 + col) <= 253868) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253869 && (row * 640 + col) <= 253874) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253875 && (row * 640 + col) <= 253880) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253881 && (row * 640 + col) <= 253883) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253884 && (row * 640 + col) <= 253889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253890 && (row * 640 + col) <= 253892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253893 && (row * 640 + col) <= 253898) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253899 && (row * 640 + col) <= 253910) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253911 && (row * 640 + col) <= 253916) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253917 && (row * 640 + col) <= 253928) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253929 && (row * 640 + col) <= 253940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253941 && (row * 640 + col) <= 253946) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253947 && (row * 640 + col) <= 253958) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253959 && (row * 640 + col) <= 253996) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 253997 && (row * 640 + col) <= 254042) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 254043 && (row * 640 + col) <= 254050) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254051 && (row * 640 + col) <= 254073) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 254074 && (row * 640 + col) <= 254231) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254232 && (row * 640 + col) <= 254234) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254235 && (row * 640 + col) <= 254268) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 254269 && (row * 640 + col) <= 254280) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 254281 && (row * 640 + col) <= 254317) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 254318 && (row * 640 + col) <= 254319) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254320 && (row * 640 + col) <= 254355) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254356 && (row * 640 + col) <= 254361) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254362 && (row * 640 + col) <= 254367) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254368 && (row * 640 + col) <= 254379) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254380 && (row * 640 + col) <= 254388) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254389 && (row * 640 + col) <= 254397) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254398 && (row * 640 + col) <= 254406) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254407 && (row * 640 + col) <= 254412) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254413 && (row * 640 + col) <= 254424) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254425 && (row * 640 + col) <= 254430) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254431 && (row * 640 + col) <= 254442) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254443 && (row * 640 + col) <= 254448) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254449 && (row * 640 + col) <= 254451) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254452 && (row * 640 + col) <= 254457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254458 && (row * 640 + col) <= 254460) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254461 && (row * 640 + col) <= 254466) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254467 && (row * 640 + col) <= 254469) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254470 && (row * 640 + col) <= 254478) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254479 && (row * 640 + col) <= 254484) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254485 && (row * 640 + col) <= 254490) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254491 && (row * 640 + col) <= 254496) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254497 && (row * 640 + col) <= 254508) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254509 && (row * 640 + col) <= 254514) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254515 && (row * 640 + col) <= 254520) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254521 && (row * 640 + col) <= 254523) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254524 && (row * 640 + col) <= 254529) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254530 && (row * 640 + col) <= 254532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254533 && (row * 640 + col) <= 254538) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254539 && (row * 640 + col) <= 254550) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254551 && (row * 640 + col) <= 254556) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254557 && (row * 640 + col) <= 254568) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254569 && (row * 640 + col) <= 254580) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254581 && (row * 640 + col) <= 254586) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254587 && (row * 640 + col) <= 254598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254599 && (row * 640 + col) <= 254636) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254637 && (row * 640 + col) <= 254682) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 254683 && (row * 640 + col) <= 254690) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254691 && (row * 640 + col) <= 254713) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 254714 && (row * 640 + col) <= 254871) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254872 && (row * 640 + col) <= 254873) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254874 && (row * 640 + col) <= 254908) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 254909 && (row * 640 + col) <= 254920) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 254921 && (row * 640 + col) <= 254957) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 254958 && (row * 640 + col) <= 254959) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254960 && (row * 640 + col) <= 254995) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 254996 && (row * 640 + col) <= 255001) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255002 && (row * 640 + col) <= 255007) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255008 && (row * 640 + col) <= 255013) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255014 && (row * 640 + col) <= 255034) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255035 && (row * 640 + col) <= 255040) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255041 && (row * 640 + col) <= 255046) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255047 && (row * 640 + col) <= 255052) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255053 && (row * 640 + col) <= 255064) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255065 && (row * 640 + col) <= 255070) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255071 && (row * 640 + col) <= 255082) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255083 && (row * 640 + col) <= 255088) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255089 && (row * 640 + col) <= 255091) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255092 && (row * 640 + col) <= 255097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255098 && (row * 640 + col) <= 255100) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255101 && (row * 640 + col) <= 255106) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255107 && (row * 640 + col) <= 255112) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255113 && (row * 640 + col) <= 255118) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255119 && (row * 640 + col) <= 255124) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255125 && (row * 640 + col) <= 255130) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255131 && (row * 640 + col) <= 255136) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255137 && (row * 640 + col) <= 255142) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255143 && (row * 640 + col) <= 255145) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255146 && (row * 640 + col) <= 255151) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255152 && (row * 640 + col) <= 255154) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255155 && (row * 640 + col) <= 255160) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255161 && (row * 640 + col) <= 255163) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255164 && (row * 640 + col) <= 255169) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255170 && (row * 640 + col) <= 255172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255173 && (row * 640 + col) <= 255178) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255179 && (row * 640 + col) <= 255190) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255191 && (row * 640 + col) <= 255196) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255197 && (row * 640 + col) <= 255208) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255209 && (row * 640 + col) <= 255214) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255215 && (row * 640 + col) <= 255226) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255227 && (row * 640 + col) <= 255232) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255233 && (row * 640 + col) <= 255235) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255236 && (row * 640 + col) <= 255241) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255242 && (row * 640 + col) <= 255276) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255277 && (row * 640 + col) <= 255322) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 255323 && (row * 640 + col) <= 255330) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255331 && (row * 640 + col) <= 255353) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 255354 && (row * 640 + col) <= 255510) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255511 && (row * 640 + col) <= 255513) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255514 && (row * 640 + col) <= 255551) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 255552 && (row * 640 + col) <= 255557) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 255558 && (row * 640 + col) <= 255597) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 255598 && (row * 640 + col) <= 255599) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255600 && (row * 640 + col) <= 255635) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255636 && (row * 640 + col) <= 255641) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255642 && (row * 640 + col) <= 255647) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255648 && (row * 640 + col) <= 255653) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255654 && (row * 640 + col) <= 255674) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255675 && (row * 640 + col) <= 255680) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255681 && (row * 640 + col) <= 255686) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255687 && (row * 640 + col) <= 255692) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255693 && (row * 640 + col) <= 255704) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255705 && (row * 640 + col) <= 255710) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255711 && (row * 640 + col) <= 255722) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255723 && (row * 640 + col) <= 255728) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255729 && (row * 640 + col) <= 255731) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255732 && (row * 640 + col) <= 255737) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255738 && (row * 640 + col) <= 255740) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255741 && (row * 640 + col) <= 255746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255747 && (row * 640 + col) <= 255752) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255753 && (row * 640 + col) <= 255758) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255759 && (row * 640 + col) <= 255764) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255765 && (row * 640 + col) <= 255770) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255771 && (row * 640 + col) <= 255776) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255777 && (row * 640 + col) <= 255782) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255783 && (row * 640 + col) <= 255785) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255786 && (row * 640 + col) <= 255791) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255792 && (row * 640 + col) <= 255794) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255795 && (row * 640 + col) <= 255800) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255801 && (row * 640 + col) <= 255803) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255804 && (row * 640 + col) <= 255809) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255810 && (row * 640 + col) <= 255812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255813 && (row * 640 + col) <= 255818) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255819 && (row * 640 + col) <= 255830) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255831 && (row * 640 + col) <= 255836) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255837 && (row * 640 + col) <= 255848) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255849 && (row * 640 + col) <= 255854) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255855 && (row * 640 + col) <= 255866) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255867 && (row * 640 + col) <= 255872) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255873 && (row * 640 + col) <= 255875) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255876 && (row * 640 + col) <= 255881) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255882 && (row * 640 + col) <= 255916) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255917 && (row * 640 + col) <= 255939) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 255940 && (row * 640 + col) <= 255944) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255945 && (row * 640 + col) <= 255962) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 255963 && (row * 640 + col) <= 255970) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 255971 && (row * 640 + col) <= 255993) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 255994 && (row * 640 + col) <= 256150) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256151 && (row * 640 + col) <= 256152) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256153 && (row * 640 + col) <= 256191) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 256192 && (row * 640 + col) <= 256197) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 256198 && (row * 640 + col) <= 256237) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 256238 && (row * 640 + col) <= 256239) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256240 && (row * 640 + col) <= 256275) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256276 && (row * 640 + col) <= 256281) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256282 && (row * 640 + col) <= 256287) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256288 && (row * 640 + col) <= 256293) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256294 && (row * 640 + col) <= 256314) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256315 && (row * 640 + col) <= 256320) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256321 && (row * 640 + col) <= 256326) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256327 && (row * 640 + col) <= 256332) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256333 && (row * 640 + col) <= 256344) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256345 && (row * 640 + col) <= 256350) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256351 && (row * 640 + col) <= 256362) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256363 && (row * 640 + col) <= 256368) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256369 && (row * 640 + col) <= 256371) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256372 && (row * 640 + col) <= 256377) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256378 && (row * 640 + col) <= 256380) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256381 && (row * 640 + col) <= 256386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256387 && (row * 640 + col) <= 256392) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256393 && (row * 640 + col) <= 256398) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256399 && (row * 640 + col) <= 256404) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256405 && (row * 640 + col) <= 256410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256411 && (row * 640 + col) <= 256416) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256417 && (row * 640 + col) <= 256422) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256423 && (row * 640 + col) <= 256425) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256426 && (row * 640 + col) <= 256431) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256432 && (row * 640 + col) <= 256434) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256435 && (row * 640 + col) <= 256440) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256441 && (row * 640 + col) <= 256443) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256444 && (row * 640 + col) <= 256449) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256450 && (row * 640 + col) <= 256452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256453 && (row * 640 + col) <= 256458) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256459 && (row * 640 + col) <= 256470) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256471 && (row * 640 + col) <= 256476) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256477 && (row * 640 + col) <= 256488) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256489 && (row * 640 + col) <= 256494) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256495 && (row * 640 + col) <= 256506) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256507 && (row * 640 + col) <= 256512) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256513 && (row * 640 + col) <= 256515) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256516 && (row * 640 + col) <= 256521) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256522 && (row * 640 + col) <= 256556) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256557 && (row * 640 + col) <= 256579) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 256580 && (row * 640 + col) <= 256584) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256585 && (row * 640 + col) <= 256602) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 256603 && (row * 640 + col) <= 256610) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256611 && (row * 640 + col) <= 256633) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 256634 && (row * 640 + col) <= 256790) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256791 && (row * 640 + col) <= 256792) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256793 && (row * 640 + col) <= 256831) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 256832 && (row * 640 + col) <= 256837) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 256838 && (row * 640 + col) <= 256877) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 256878 && (row * 640 + col) <= 256879) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256880 && (row * 640 + col) <= 256915) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256916 && (row * 640 + col) <= 256921) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256922 && (row * 640 + col) <= 256927) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256928 && (row * 640 + col) <= 256933) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256934 && (row * 640 + col) <= 256954) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256955 && (row * 640 + col) <= 256960) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256961 && (row * 640 + col) <= 256966) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256967 && (row * 640 + col) <= 256972) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256973 && (row * 640 + col) <= 256984) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 256985 && (row * 640 + col) <= 256990) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256991 && (row * 640 + col) <= 257002) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257003 && (row * 640 + col) <= 257008) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257009 && (row * 640 + col) <= 257011) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257012 && (row * 640 + col) <= 257017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257018 && (row * 640 + col) <= 257020) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257021 && (row * 640 + col) <= 257026) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257027 && (row * 640 + col) <= 257032) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257033 && (row * 640 + col) <= 257038) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257039 && (row * 640 + col) <= 257044) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257045 && (row * 640 + col) <= 257050) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257051 && (row * 640 + col) <= 257056) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257057 && (row * 640 + col) <= 257062) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257063 && (row * 640 + col) <= 257065) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257066 && (row * 640 + col) <= 257071) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257072 && (row * 640 + col) <= 257074) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257075 && (row * 640 + col) <= 257080) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257081 && (row * 640 + col) <= 257083) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257084 && (row * 640 + col) <= 257089) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257090 && (row * 640 + col) <= 257092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257093 && (row * 640 + col) <= 257098) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257099 && (row * 640 + col) <= 257110) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257111 && (row * 640 + col) <= 257116) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257117 && (row * 640 + col) <= 257128) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257129 && (row * 640 + col) <= 257134) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257135 && (row * 640 + col) <= 257146) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257147 && (row * 640 + col) <= 257152) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257153 && (row * 640 + col) <= 257155) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257156 && (row * 640 + col) <= 257161) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257162 && (row * 640 + col) <= 257196) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257197 && (row * 640 + col) <= 257219) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 257220 && (row * 640 + col) <= 257224) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257225 && (row * 640 + col) <= 257239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 257240 && (row * 640 + col) <= 257429) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257430 && (row * 640 + col) <= 257432) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257433 && (row * 640 + col) <= 257471) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 257472 && (row * 640 + col) <= 257477) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 257478 && (row * 640 + col) <= 257517) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 257518 && (row * 640 + col) <= 257518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257519 && (row * 640 + col) <= 257555) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257556 && (row * 640 + col) <= 257561) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257562 && (row * 640 + col) <= 257567) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257568 && (row * 640 + col) <= 257573) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257574 && (row * 640 + col) <= 257594) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257595 && (row * 640 + col) <= 257600) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257601 && (row * 640 + col) <= 257606) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257607 && (row * 640 + col) <= 257612) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257613 && (row * 640 + col) <= 257624) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257625 && (row * 640 + col) <= 257630) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257631 && (row * 640 + col) <= 257642) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257643 && (row * 640 + col) <= 257648) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257649 && (row * 640 + col) <= 257651) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257652 && (row * 640 + col) <= 257657) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257658 && (row * 640 + col) <= 257660) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257661 && (row * 640 + col) <= 257666) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257667 && (row * 640 + col) <= 257672) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257673 && (row * 640 + col) <= 257678) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257679 && (row * 640 + col) <= 257684) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257685 && (row * 640 + col) <= 257690) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257691 && (row * 640 + col) <= 257696) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257697 && (row * 640 + col) <= 257702) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257703 && (row * 640 + col) <= 257705) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257706 && (row * 640 + col) <= 257711) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257712 && (row * 640 + col) <= 257714) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257715 && (row * 640 + col) <= 257720) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257721 && (row * 640 + col) <= 257723) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257724 && (row * 640 + col) <= 257729) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257730 && (row * 640 + col) <= 257732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257733 && (row * 640 + col) <= 257738) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257739 && (row * 640 + col) <= 257750) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257751 && (row * 640 + col) <= 257756) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257757 && (row * 640 + col) <= 257768) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257769 && (row * 640 + col) <= 257774) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257775 && (row * 640 + col) <= 257786) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257787 && (row * 640 + col) <= 257792) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257793 && (row * 640 + col) <= 257795) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257796 && (row * 640 + col) <= 257801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257802 && (row * 640 + col) <= 257836) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257837 && (row * 640 + col) <= 257859) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 257860 && (row * 640 + col) <= 257864) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 257865 && (row * 640 + col) <= 257879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 257880 && (row * 640 + col) <= 258069) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258070 && (row * 640 + col) <= 258071) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258072 && (row * 640 + col) <= 258111) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 258112 && (row * 640 + col) <= 258117) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 258118 && (row * 640 + col) <= 258156) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 258157 && (row * 640 + col) <= 258158) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258159 && (row * 640 + col) <= 258169) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258170 && (row * 640 + col) <= 258173) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258174 && (row * 640 + col) <= 258195) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258196 && (row * 640 + col) <= 258201) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258202 && (row * 640 + col) <= 258207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258208 && (row * 640 + col) <= 258213) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258214 && (row * 640 + col) <= 258234) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258235 && (row * 640 + col) <= 258240) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258241 && (row * 640 + col) <= 258246) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258247 && (row * 640 + col) <= 258252) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258253 && (row * 640 + col) <= 258264) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258265 && (row * 640 + col) <= 258270) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258271 && (row * 640 + col) <= 258282) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258283 && (row * 640 + col) <= 258288) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258289 && (row * 640 + col) <= 258291) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258292 && (row * 640 + col) <= 258297) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258298 && (row * 640 + col) <= 258300) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258301 && (row * 640 + col) <= 258306) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258307 && (row * 640 + col) <= 258312) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258313 && (row * 640 + col) <= 258318) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258319 && (row * 640 + col) <= 258324) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258325 && (row * 640 + col) <= 258330) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258331 && (row * 640 + col) <= 258336) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258337 && (row * 640 + col) <= 258342) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258343 && (row * 640 + col) <= 258345) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258346 && (row * 640 + col) <= 258351) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258352 && (row * 640 + col) <= 258354) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258355 && (row * 640 + col) <= 258360) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258361 && (row * 640 + col) <= 258363) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258364 && (row * 640 + col) <= 258369) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258370 && (row * 640 + col) <= 258372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258373 && (row * 640 + col) <= 258378) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258379 && (row * 640 + col) <= 258390) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258391 && (row * 640 + col) <= 258396) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258397 && (row * 640 + col) <= 258408) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258409 && (row * 640 + col) <= 258414) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258415 && (row * 640 + col) <= 258426) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258427 && (row * 640 + col) <= 258432) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258433 && (row * 640 + col) <= 258435) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258436 && (row * 640 + col) <= 258441) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258442 && (row * 640 + col) <= 258476) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258477 && (row * 640 + col) <= 258499) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 258500 && (row * 640 + col) <= 258504) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258505 && (row * 640 + col) <= 258519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 258520 && (row * 640 + col) <= 258709) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258710 && (row * 640 + col) <= 258711) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258712 && (row * 640 + col) <= 258751) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 258752 && (row * 640 + col) <= 258757) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 258758 && (row * 640 + col) <= 258796) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 258797 && (row * 640 + col) <= 258798) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258799 && (row * 640 + col) <= 258809) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258810 && (row * 640 + col) <= 258813) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258814 && (row * 640 + col) <= 258835) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258836 && (row * 640 + col) <= 258841) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258842 && (row * 640 + col) <= 258847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258848 && (row * 640 + col) <= 258853) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258854 && (row * 640 + col) <= 258856) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258857 && (row * 640 + col) <= 258862) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258863 && (row * 640 + col) <= 258865) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258866 && (row * 640 + col) <= 258871) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258872 && (row * 640 + col) <= 258874) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258875 && (row * 640 + col) <= 258880) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258881 && (row * 640 + col) <= 258886) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258887 && (row * 640 + col) <= 258892) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258893 && (row * 640 + col) <= 258904) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258905 && (row * 640 + col) <= 258910) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258911 && (row * 640 + col) <= 258913) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258914 && (row * 640 + col) <= 258919) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258920 && (row * 640 + col) <= 258922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258923 && (row * 640 + col) <= 258928) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258929 && (row * 640 + col) <= 258931) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258932 && (row * 640 + col) <= 258937) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258938 && (row * 640 + col) <= 258940) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258941 && (row * 640 + col) <= 258946) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258947 && (row * 640 + col) <= 258952) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258953 && (row * 640 + col) <= 258958) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258959 && (row * 640 + col) <= 258964) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258965 && (row * 640 + col) <= 258970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258971 && (row * 640 + col) <= 258976) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258977 && (row * 640 + col) <= 258982) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258983 && (row * 640 + col) <= 258985) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258986 && (row * 640 + col) <= 258991) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258992 && (row * 640 + col) <= 258994) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 258995 && (row * 640 + col) <= 259000) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259001 && (row * 640 + col) <= 259003) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259004 && (row * 640 + col) <= 259009) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259010 && (row * 640 + col) <= 259012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259013 && (row * 640 + col) <= 259018) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259019 && (row * 640 + col) <= 259030) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259031 && (row * 640 + col) <= 259036) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259037 && (row * 640 + col) <= 259048) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259049 && (row * 640 + col) <= 259054) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259055 && (row * 640 + col) <= 259057) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259058 && (row * 640 + col) <= 259063) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259064 && (row * 640 + col) <= 259066) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259067 && (row * 640 + col) <= 259072) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259073 && (row * 640 + col) <= 259075) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259076 && (row * 640 + col) <= 259081) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259082 && (row * 640 + col) <= 259116) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259117 && (row * 640 + col) <= 259127) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 259128 && (row * 640 + col) <= 259150) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259151 && (row * 640 + col) <= 259159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 259160 && (row * 640 + col) <= 259348) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259349 && (row * 640 + col) <= 259351) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259352 && (row * 640 + col) <= 259391) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 259392 && (row * 640 + col) <= 259397) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 259398 && (row * 640 + col) <= 259435) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 259436 && (row * 640 + col) <= 259437) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259438 && (row * 640 + col) <= 259449) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259450 && (row * 640 + col) <= 259453) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259454 && (row * 640 + col) <= 259475) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259476 && (row * 640 + col) <= 259481) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259482 && (row * 640 + col) <= 259487) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259488 && (row * 640 + col) <= 259493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259494 && (row * 640 + col) <= 259496) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259497 && (row * 640 + col) <= 259502) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259503 && (row * 640 + col) <= 259505) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259506 && (row * 640 + col) <= 259511) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259512 && (row * 640 + col) <= 259514) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259515 && (row * 640 + col) <= 259520) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259521 && (row * 640 + col) <= 259526) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259527 && (row * 640 + col) <= 259532) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259533 && (row * 640 + col) <= 259544) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259545 && (row * 640 + col) <= 259550) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259551 && (row * 640 + col) <= 259553) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259554 && (row * 640 + col) <= 259559) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259560 && (row * 640 + col) <= 259562) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259563 && (row * 640 + col) <= 259568) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259569 && (row * 640 + col) <= 259571) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259572 && (row * 640 + col) <= 259577) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259578 && (row * 640 + col) <= 259580) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259581 && (row * 640 + col) <= 259586) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259587 && (row * 640 + col) <= 259592) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259593 && (row * 640 + col) <= 259598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259599 && (row * 640 + col) <= 259604) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259605 && (row * 640 + col) <= 259610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259611 && (row * 640 + col) <= 259616) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259617 && (row * 640 + col) <= 259622) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259623 && (row * 640 + col) <= 259625) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259626 && (row * 640 + col) <= 259631) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259632 && (row * 640 + col) <= 259634) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259635 && (row * 640 + col) <= 259640) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259641 && (row * 640 + col) <= 259643) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259644 && (row * 640 + col) <= 259649) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259650 && (row * 640 + col) <= 259652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259653 && (row * 640 + col) <= 259658) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259659 && (row * 640 + col) <= 259670) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259671 && (row * 640 + col) <= 259676) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259677 && (row * 640 + col) <= 259688) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259689 && (row * 640 + col) <= 259694) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259695 && (row * 640 + col) <= 259697) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259698 && (row * 640 + col) <= 259703) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259704 && (row * 640 + col) <= 259706) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259707 && (row * 640 + col) <= 259712) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259713 && (row * 640 + col) <= 259715) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259716 && (row * 640 + col) <= 259721) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259722 && (row * 640 + col) <= 259756) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259757 && (row * 640 + col) <= 259767) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 259768 && (row * 640 + col) <= 259790) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259791 && (row * 640 + col) <= 259799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 259800 && (row * 640 + col) <= 259988) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 259989 && (row * 640 + col) <= 259990) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259991 && (row * 640 + col) <= 260031) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 260032 && (row * 640 + col) <= 260037) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 260038 && (row * 640 + col) <= 260075) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 260076 && (row * 640 + col) <= 260077) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260078 && (row * 640 + col) <= 260089) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260090 && (row * 640 + col) <= 260093) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260094 && (row * 640 + col) <= 260115) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260116 && (row * 640 + col) <= 260121) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260122 && (row * 640 + col) <= 260127) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260128 && (row * 640 + col) <= 260133) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260134 && (row * 640 + col) <= 260136) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260137 && (row * 640 + col) <= 260142) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260143 && (row * 640 + col) <= 260145) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260146 && (row * 640 + col) <= 260151) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260152 && (row * 640 + col) <= 260154) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260155 && (row * 640 + col) <= 260160) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260161 && (row * 640 + col) <= 260166) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260167 && (row * 640 + col) <= 260172) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260173 && (row * 640 + col) <= 260184) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260185 && (row * 640 + col) <= 260190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260191 && (row * 640 + col) <= 260193) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260194 && (row * 640 + col) <= 260199) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260200 && (row * 640 + col) <= 260202) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260203 && (row * 640 + col) <= 260208) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260209 && (row * 640 + col) <= 260211) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260212 && (row * 640 + col) <= 260217) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260218 && (row * 640 + col) <= 260220) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260221 && (row * 640 + col) <= 260226) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260227 && (row * 640 + col) <= 260232) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260233 && (row * 640 + col) <= 260238) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260239 && (row * 640 + col) <= 260244) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260245 && (row * 640 + col) <= 260250) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260251 && (row * 640 + col) <= 260256) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260257 && (row * 640 + col) <= 260262) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260263 && (row * 640 + col) <= 260265) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260266 && (row * 640 + col) <= 260271) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260272 && (row * 640 + col) <= 260274) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260275 && (row * 640 + col) <= 260280) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260281 && (row * 640 + col) <= 260283) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260284 && (row * 640 + col) <= 260289) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260290 && (row * 640 + col) <= 260292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260293 && (row * 640 + col) <= 260298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260299 && (row * 640 + col) <= 260310) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260311 && (row * 640 + col) <= 260316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260317 && (row * 640 + col) <= 260328) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260329 && (row * 640 + col) <= 260334) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260335 && (row * 640 + col) <= 260337) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260338 && (row * 640 + col) <= 260343) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260344 && (row * 640 + col) <= 260346) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260347 && (row * 640 + col) <= 260352) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260353 && (row * 640 + col) <= 260355) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260356 && (row * 640 + col) <= 260361) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260362 && (row * 640 + col) <= 260396) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260397 && (row * 640 + col) <= 260407) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 260408 && (row * 640 + col) <= 260430) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260431 && (row * 640 + col) <= 260439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 260440 && (row * 640 + col) <= 260628) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260629 && (row * 640 + col) <= 260630) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260631 && (row * 640 + col) <= 260671) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 260672 && (row * 640 + col) <= 260677) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 260678 && (row * 640 + col) <= 260714) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 260715 && (row * 640 + col) <= 260717) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260718 && (row * 640 + col) <= 260755) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260756 && (row * 640 + col) <= 260761) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260762 && (row * 640 + col) <= 260767) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260768 && (row * 640 + col) <= 260782) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260783 && (row * 640 + col) <= 260785) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260786 && (row * 640 + col) <= 260800) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260801 && (row * 640 + col) <= 260806) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260807 && (row * 640 + col) <= 260812) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260813 && (row * 640 + col) <= 260824) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260825 && (row * 640 + col) <= 260839) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260840 && (row * 640 + col) <= 260842) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260843 && (row * 640 + col) <= 260857) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260858 && (row * 640 + col) <= 260860) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260861 && (row * 640 + col) <= 260866) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260867 && (row * 640 + col) <= 260872) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260873 && (row * 640 + col) <= 260878) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260879 && (row * 640 + col) <= 260884) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260885 && (row * 640 + col) <= 260890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260891 && (row * 640 + col) <= 260896) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260897 && (row * 640 + col) <= 260902) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260903 && (row * 640 + col) <= 260905) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260906 && (row * 640 + col) <= 260911) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260912 && (row * 640 + col) <= 260914) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260915 && (row * 640 + col) <= 260929) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260930 && (row * 640 + col) <= 260932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260933 && (row * 640 + col) <= 260947) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260948 && (row * 640 + col) <= 260950) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260951 && (row * 640 + col) <= 260965) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260966 && (row * 640 + col) <= 260968) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260969 && (row * 640 + col) <= 260983) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260984 && (row * 640 + col) <= 260986) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260987 && (row * 640 + col) <= 260992) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260993 && (row * 640 + col) <= 260995) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 260996 && (row * 640 + col) <= 261001) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261002 && (row * 640 + col) <= 261036) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261037 && (row * 640 + col) <= 261047) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 261048 && (row * 640 + col) <= 261070) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261071 && (row * 640 + col) <= 261079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 261080 && (row * 640 + col) <= 261268) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261269 && (row * 640 + col) <= 261270) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261271 && (row * 640 + col) <= 261311) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 261312 && (row * 640 + col) <= 261317) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 261318 && (row * 640 + col) <= 261353) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 261354 && (row * 640 + col) <= 261356) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261357 && (row * 640 + col) <= 261395) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261396 && (row * 640 + col) <= 261401) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261402 && (row * 640 + col) <= 261407) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261408 && (row * 640 + col) <= 261422) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261423 && (row * 640 + col) <= 261425) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261426 && (row * 640 + col) <= 261440) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261441 && (row * 640 + col) <= 261446) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261447 && (row * 640 + col) <= 261452) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261453 && (row * 640 + col) <= 261464) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261465 && (row * 640 + col) <= 261479) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261480 && (row * 640 + col) <= 261482) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261483 && (row * 640 + col) <= 261497) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261498 && (row * 640 + col) <= 261500) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261501 && (row * 640 + col) <= 261506) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261507 && (row * 640 + col) <= 261512) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261513 && (row * 640 + col) <= 261518) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261519 && (row * 640 + col) <= 261524) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261525 && (row * 640 + col) <= 261530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261531 && (row * 640 + col) <= 261536) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261537 && (row * 640 + col) <= 261542) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261543 && (row * 640 + col) <= 261545) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261546 && (row * 640 + col) <= 261551) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261552 && (row * 640 + col) <= 261554) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261555 && (row * 640 + col) <= 261569) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261570 && (row * 640 + col) <= 261572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261573 && (row * 640 + col) <= 261587) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261588 && (row * 640 + col) <= 261590) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261591 && (row * 640 + col) <= 261605) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261606 && (row * 640 + col) <= 261608) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261609 && (row * 640 + col) <= 261623) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261624 && (row * 640 + col) <= 261626) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261627 && (row * 640 + col) <= 261632) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261633 && (row * 640 + col) <= 261635) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261636 && (row * 640 + col) <= 261641) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261642 && (row * 640 + col) <= 261676) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261677 && (row * 640 + col) <= 261687) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 261688 && (row * 640 + col) <= 261710) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261711 && (row * 640 + col) <= 261719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 261720 && (row * 640 + col) <= 261908) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 261909 && (row * 640 + col) <= 261910) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261911 && (row * 640 + col) <= 261951) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 261952 && (row * 640 + col) <= 261957) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 261958 && (row * 640 + col) <= 261992) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 261993 && (row * 640 + col) <= 261995) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261996 && (row * 640 + col) <= 262035) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262036 && (row * 640 + col) <= 262041) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262042 && (row * 640 + col) <= 262047) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262048 && (row * 640 + col) <= 262062) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262063 && (row * 640 + col) <= 262065) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262066 && (row * 640 + col) <= 262080) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262081 && (row * 640 + col) <= 262086) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262087 && (row * 640 + col) <= 262092) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262093 && (row * 640 + col) <= 262104) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262105 && (row * 640 + col) <= 262119) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262120 && (row * 640 + col) <= 262122) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262123 && (row * 640 + col) <= 262137) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262138 && (row * 640 + col) <= 262140) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262141 && (row * 640 + col) <= 262146) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262147 && (row * 640 + col) <= 262152) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262153 && (row * 640 + col) <= 262158) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262159 && (row * 640 + col) <= 262164) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262165 && (row * 640 + col) <= 262170) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262171 && (row * 640 + col) <= 262176) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262177 && (row * 640 + col) <= 262182) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262183 && (row * 640 + col) <= 262185) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262186 && (row * 640 + col) <= 262191) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262192 && (row * 640 + col) <= 262194) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262195 && (row * 640 + col) <= 262209) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262210 && (row * 640 + col) <= 262212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262213 && (row * 640 + col) <= 262227) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262228 && (row * 640 + col) <= 262230) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262231 && (row * 640 + col) <= 262245) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262246 && (row * 640 + col) <= 262248) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262249 && (row * 640 + col) <= 262263) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262264 && (row * 640 + col) <= 262266) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262267 && (row * 640 + col) <= 262272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262273 && (row * 640 + col) <= 262275) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262276 && (row * 640 + col) <= 262281) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262282 && (row * 640 + col) <= 262316) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262317 && (row * 640 + col) <= 262327) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 262328 && (row * 640 + col) <= 262350) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262351 && (row * 640 + col) <= 262359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 262360 && (row * 640 + col) <= 262548) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262549 && (row * 640 + col) <= 262550) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262551 && (row * 640 + col) <= 262591) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 262592 && (row * 640 + col) <= 262597) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 262598 && (row * 640 + col) <= 262631) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 262632 && (row * 640 + col) <= 262634) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262635 && (row * 640 + col) <= 262990) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 262991 && (row * 640 + col) <= 262999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 263000 && (row * 640 + col) <= 263188) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 263189 && (row * 640 + col) <= 263190) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263191 && (row * 640 + col) <= 263270) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 263271 && (row * 640 + col) <= 263274) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263275 && (row * 640 + col) <= 263630) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 263631 && (row * 640 + col) <= 263639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 263640 && (row * 640 + col) <= 263828) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 263829 && (row * 640 + col) <= 263830) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263831 && (row * 640 + col) <= 263908) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 263909 && (row * 640 + col) <= 263912) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263913 && (row * 640 + col) <= 264270) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 264271 && (row * 640 + col) <= 264279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 264280 && (row * 640 + col) <= 264468) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 264469 && (row * 640 + col) <= 264471) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264472 && (row * 640 + col) <= 264546) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 264547 && (row * 640 + col) <= 264551) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264552 && (row * 640 + col) <= 264910) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 264911 && (row * 640 + col) <= 264919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 264920 && (row * 640 + col) <= 265109) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 265110 && (row * 640 + col) <= 265111) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265112 && (row * 640 + col) <= 265184) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 265185 && (row * 640 + col) <= 265189) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265190 && (row * 640 + col) <= 265550) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 265551 && (row * 640 + col) <= 265559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 265560 && (row * 640 + col) <= 265749) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 265750 && (row * 640 + col) <= 265751) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265752 && (row * 640 + col) <= 265809) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 265810 && (row * 640 + col) <= 265827) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265828 && (row * 640 + col) <= 266190) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 266191 && (row * 640 + col) <= 266199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 266200 && (row * 640 + col) <= 266389) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 266390 && (row * 640 + col) <= 266392) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 266393 && (row * 640 + col) <= 266437) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 266438 && (row * 640 + col) <= 266465) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 266466 && (row * 640 + col) <= 267030) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 267031 && (row * 640 + col) <= 267032) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 267033 && (row * 640 + col) <= 267071) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 267072 && (row * 640 + col) <= 267090) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 267091 && (row * 640 + col) <= 267670) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 267671 && (row * 640 + col) <= 267673) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 267674 && (row * 640 + col) <= 267708) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 267709 && (row * 640 + col) <= 267718) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 267719 && (row * 640 + col) <= 268311) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 268312 && (row * 640 + col) <= 268314) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 268315 && (row * 640 + col) <= 268345) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 268346 && (row * 640 + col) <= 268352) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 268353 && (row * 640 + col) <= 268951) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 268952 && (row * 640 + col) <= 268954) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 268955 && (row * 640 + col) <= 268983) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 268984 && (row * 640 + col) <= 268989) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 268990 && (row * 640 + col) <= 269592) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 269593 && (row * 640 + col) <= 269595) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 269596 && (row * 640 + col) <= 269621) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 269622 && (row * 640 + col) <= 269626) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 269627 && (row * 640 + col) <= 270233) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 270234 && (row * 640 + col) <= 270236) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 270237 && (row * 640 + col) <= 270259) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 270260 && (row * 640 + col) <= 270264) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 270265 && (row * 640 + col) <= 270874) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 270875 && (row * 640 + col) <= 270877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 270878 && (row * 640 + col) <= 270896) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 270897 && (row * 640 + col) <= 270902) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 270903 && (row * 640 + col) <= 271515) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 271516 && (row * 640 + col) <= 271519) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 271520 && (row * 640 + col) <= 271534) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 271535 && (row * 640 + col) <= 271540) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 271541 && (row * 640 + col) <= 272156) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 272157 && (row * 640 + col) <= 272162) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 272163 && (row * 640 + col) <= 272170) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 272171 && (row * 640 + col) <= 272177) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 272178 && (row * 640 + col) <= 272798) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 272799 && (row * 640 + col) <= 272815) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 272816 && (row * 640 + col) <= 273441) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 273442 && (row * 640 + col) <= 273451) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 273452 && (row * 640 + col) <= 284159) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 284160 && (row * 640 + col) < 307200) color_data <= 12'b010010000001; else
        color_data <= 12'b000000000000;
    end
endmodule
