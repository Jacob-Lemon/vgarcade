module seven_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "distributed" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		10'b0000100100: color_data = 12'b000000000000;
		10'b0000100101: color_data = 12'b000000000000;
		10'b0000100110: color_data = 12'b000000000000;
		10'b0000100111: color_data = 12'b000000000000;
		10'b0000101000: color_data = 12'b000000000000;
		10'b0000101001: color_data = 12'b000000000000;
		10'b0000101010: color_data = 12'b000000000000;
		10'b0000101011: color_data = 12'b000000000000;
		10'b0000101100: color_data = 12'b000000000000;
		10'b0000101101: color_data = 12'b000000000000;
		10'b0000101110: color_data = 12'b000000000000;
		10'b0000101111: color_data = 12'b000000000000;
		10'b0000110000: color_data = 12'b000000000000;
		10'b0000110001: color_data = 12'b000000000000;
		10'b0000110010: color_data = 12'b000000000000;
		10'b0000110011: color_data = 12'b000000000000;
		10'b0001000010: color_data = 12'b000000000000;
		10'b0001000011: color_data = 12'b000000000000;
		10'b0001000100: color_data = 12'b000000000000;
		10'b0001000101: color_data = 12'b000000000000;
		10'b0001000110: color_data = 12'b000000000000;
		10'b0001000111: color_data = 12'b000000000000;
		10'b0001001000: color_data = 12'b000000000000;
		10'b0001001001: color_data = 12'b000000000000;
		10'b0001001010: color_data = 12'b000000000000;
		10'b0001001011: color_data = 12'b000000000000;
		10'b0001001100: color_data = 12'b000000000000;
		10'b0001001101: color_data = 12'b000000000000;
		10'b0001001110: color_data = 12'b000000000000;
		10'b0001001111: color_data = 12'b000000000000;
		10'b0001010000: color_data = 12'b000000000000;
		10'b0001010001: color_data = 12'b000000000000;
		10'b0001010010: color_data = 12'b000000000000;
		10'b0001010011: color_data = 12'b000000000000;
		10'b0001010100: color_data = 12'b000000000000;
		10'b0001010101: color_data = 12'b000000000000;
		10'b0001100010: color_data = 12'b000000000000;
		10'b0001100011: color_data = 12'b000000000000;
		10'b0001100100: color_data = 12'b000000000000;
		10'b0001100101: color_data = 12'b000000000000;
		10'b0001100110: color_data = 12'b000000000000;
		10'b0001100111: color_data = 12'b000000000000;
		10'b0001101000: color_data = 12'b000000000000;
		10'b0001101001: color_data = 12'b000000000000;
		10'b0001101010: color_data = 12'b000000000000;
		10'b0001101011: color_data = 12'b000000000000;
		10'b0001101100: color_data = 12'b000000000000;
		10'b0001101101: color_data = 12'b000000000000;
		10'b0001101110: color_data = 12'b000000000000;
		10'b0001101111: color_data = 12'b000000000000;
		10'b0001110000: color_data = 12'b000000000000;
		10'b0001110001: color_data = 12'b000000000000;
		10'b0001110010: color_data = 12'b000000000000;
		10'b0001110011: color_data = 12'b000000000000;
		10'b0001110100: color_data = 12'b000000000000;
		10'b0001110101: color_data = 12'b000000000000;
		10'b0001110110: color_data = 12'b000000000000;
		10'b0010000010: color_data = 12'b000000000000;
		10'b0010000011: color_data = 12'b000000000000;
		10'b0010000100: color_data = 12'b000000000000;
		10'b0010000101: color_data = 12'b000000000000;
		10'b0010000110: color_data = 12'b000000000000;
		10'b0010000111: color_data = 12'b000000000000;
		10'b0010001000: color_data = 12'b000000000000;
		10'b0010001001: color_data = 12'b000000000000;
		10'b0010001010: color_data = 12'b000000000000;
		10'b0010001011: color_data = 12'b000000000000;
		10'b0010001100: color_data = 12'b000000000000;
		10'b0010001101: color_data = 12'b000000000000;
		10'b0010001110: color_data = 12'b000000000000;
		10'b0010001111: color_data = 12'b000000000000;
		10'b0010010000: color_data = 12'b000000000000;
		10'b0010010001: color_data = 12'b000000000000;
		10'b0010010010: color_data = 12'b000000000000;
		10'b0010010011: color_data = 12'b000000000000;
		10'b0010010100: color_data = 12'b000000000000;
		10'b0010010101: color_data = 12'b000000000000;
		10'b0010010110: color_data = 12'b000000000000;
		10'b0010100011: color_data = 12'b000000000000;
		10'b0010100100: color_data = 12'b000000000000;
		10'b0010100101: color_data = 12'b000000000000;
		10'b0010100110: color_data = 12'b000000000000;
		10'b0010100111: color_data = 12'b000000000000;
		10'b0010101000: color_data = 12'b000000000000;
		10'b0010101001: color_data = 12'b000000000000;
		10'b0010101010: color_data = 12'b000000000000;
		10'b0010101011: color_data = 12'b000000000000;
		10'b0010101100: color_data = 12'b000000000000;
		10'b0010101101: color_data = 12'b000000000000;
		10'b0010101110: color_data = 12'b000000000000;
		10'b0010101111: color_data = 12'b000000000000;
		10'b0010110000: color_data = 12'b000000000000;
		10'b0010110001: color_data = 12'b000000000000;
		10'b0010110010: color_data = 12'b000000000000;
		10'b0010110011: color_data = 12'b000000000000;
		10'b0010110100: color_data = 12'b000000000000;
		10'b0010110101: color_data = 12'b000000000000;
		10'b0010110110: color_data = 12'b000000000000;
		10'b0011010000: color_data = 12'b000000000000;
		10'b0011010001: color_data = 12'b000000000000;
		10'b0011010010: color_data = 12'b000000000000;
		10'b0011010011: color_data = 12'b000000000000;
		10'b0011010100: color_data = 12'b000000000000;
		10'b0011010101: color_data = 12'b000000000000;
		10'b0011101111: color_data = 12'b000000000000;
		10'b0011110000: color_data = 12'b000000000000;
		10'b0011110001: color_data = 12'b000000000000;
		10'b0011110010: color_data = 12'b000000000000;
		10'b0011110011: color_data = 12'b000000000000;
		10'b0011110100: color_data = 12'b000000000000;
		10'b0011110101: color_data = 12'b000000000000;
		10'b0100001111: color_data = 12'b000000000000;
		10'b0100010000: color_data = 12'b000000000000;
		10'b0100010001: color_data = 12'b000000000000;
		10'b0100010010: color_data = 12'b000000000000;
		10'b0100010011: color_data = 12'b000000000000;
		10'b0100010100: color_data = 12'b000000000000;
		10'b0100101110: color_data = 12'b000000000000;
		10'b0100101111: color_data = 12'b000000000000;
		10'b0100110000: color_data = 12'b000000000000;
		10'b0100110001: color_data = 12'b000000000000;
		10'b0100110010: color_data = 12'b000000000000;
		10'b0100110011: color_data = 12'b000000000000;
		10'b0101001101: color_data = 12'b000000000000;
		10'b0101001110: color_data = 12'b000000000000;
		10'b0101001111: color_data = 12'b000000000000;
		10'b0101010000: color_data = 12'b000000000000;
		10'b0101010001: color_data = 12'b000000000000;
		10'b0101010010: color_data = 12'b000000000000;
		10'b0101010011: color_data = 12'b000000000000;
		10'b0101101101: color_data = 12'b000000000000;
		10'b0101101110: color_data = 12'b000000000000;
		10'b0101101111: color_data = 12'b000000000000;
		10'b0101110000: color_data = 12'b000000000000;
		10'b0101110001: color_data = 12'b000000000000;
		10'b0101110010: color_data = 12'b000000000000;
		10'b0110001100: color_data = 12'b000000000000;
		10'b0110001101: color_data = 12'b000000000000;
		10'b0110001110: color_data = 12'b000000000000;
		10'b0110001111: color_data = 12'b000000000000;
		10'b0110010000: color_data = 12'b000000000000;
		10'b0110010001: color_data = 12'b000000000000;
		10'b0110101011: color_data = 12'b000000000000;
		10'b0110101100: color_data = 12'b000000000000;
		10'b0110101101: color_data = 12'b000000000000;
		10'b0110101110: color_data = 12'b000000000000;
		10'b0110101111: color_data = 12'b000000000000;
		10'b0110110000: color_data = 12'b000000000000;
		10'b0111001011: color_data = 12'b000000000000;
		10'b0111001100: color_data = 12'b000000000000;
		10'b0111001101: color_data = 12'b000000000000;
		10'b0111001110: color_data = 12'b000000000000;
		10'b0111001111: color_data = 12'b000000000000;
		10'b0111010000: color_data = 12'b000000000000;
		10'b0111101010: color_data = 12'b000000000000;
		10'b0111101011: color_data = 12'b000000000000;
		10'b0111101100: color_data = 12'b000000000000;
		10'b0111101101: color_data = 12'b000000000000;
		10'b0111101110: color_data = 12'b000000000000;
		10'b0111101111: color_data = 12'b000000000000;
		10'b1000001001: color_data = 12'b000000000000;
		10'b1000001010: color_data = 12'b000000000000;
		10'b1000001011: color_data = 12'b000000000000;
		10'b1000001100: color_data = 12'b000000000000;
		10'b1000001101: color_data = 12'b000000000000;
		10'b1000001110: color_data = 12'b000000000000;
		10'b1000101001: color_data = 12'b000000000000;
		10'b1000101010: color_data = 12'b000000000000;
		10'b1000101011: color_data = 12'b000000000000;
		10'b1000101100: color_data = 12'b000000000000;
		10'b1000101101: color_data = 12'b000000000000;
		10'b1000101110: color_data = 12'b000000000000;
		10'b1001001000: color_data = 12'b000000000000;
		10'b1001001001: color_data = 12'b000000000000;
		10'b1001001010: color_data = 12'b000000000000;
		10'b1001001011: color_data = 12'b000000000000;
		10'b1001001100: color_data = 12'b000000000000;
		10'b1001001101: color_data = 12'b000000000000;
		10'b1001100111: color_data = 12'b000000000000;
		10'b1001101000: color_data = 12'b000000000000;
		10'b1001101001: color_data = 12'b000000000000;
		10'b1001101010: color_data = 12'b000000000000;
		10'b1001101011: color_data = 12'b000000000000;
		10'b1001101100: color_data = 12'b000000000000;
		10'b1010000111: color_data = 12'b000000000000;
		10'b1010001000: color_data = 12'b000000000000;
		10'b1010001001: color_data = 12'b000000000000;
		10'b1010001010: color_data = 12'b000000000000;
		10'b1010001011: color_data = 12'b000000000000;
		10'b1010001100: color_data = 12'b000000000000;
		10'b1010100110: color_data = 12'b000000000000;
		10'b1010100111: color_data = 12'b000000000000;
		10'b1010101000: color_data = 12'b000000000000;
		10'b1010101001: color_data = 12'b000000000000;
		10'b1010101010: color_data = 12'b000000000000;
		10'b1010101011: color_data = 12'b000000000000;
		10'b1011000101: color_data = 12'b000000000000;
		10'b1011000110: color_data = 12'b000000000000;
		10'b1011000111: color_data = 12'b000000000000;
		10'b1011001000: color_data = 12'b000000000000;
		10'b1011001001: color_data = 12'b000000000000;
		10'b1011001010: color_data = 12'b000000000000;
		10'b1011100101: color_data = 12'b000000000000;
		10'b1011100110: color_data = 12'b000000000000;
		10'b1011100111: color_data = 12'b000000000000;
		10'b1011101000: color_data = 12'b000000000000;
		10'b1011101001: color_data = 12'b000000000000;
		10'b1011101010: color_data = 12'b000000000000;
		10'b1100000100: color_data = 12'b000000000000;
		10'b1100000101: color_data = 12'b000000000000;
		10'b1100000110: color_data = 12'b000000000000;
		10'b1100000111: color_data = 12'b000000000000;
		10'b1100001000: color_data = 12'b000000000000;
		10'b1100001001: color_data = 12'b000000000000;
		10'b1100100011: color_data = 12'b000000000000;
		10'b1100100100: color_data = 12'b000000000000;
		10'b1100100101: color_data = 12'b000000000000;
		10'b1100100110: color_data = 12'b000000000000;
		10'b1100100111: color_data = 12'b000000000000;
		10'b1100101000: color_data = 12'b000000000000;
		10'b1101000011: color_data = 12'b000000000000;
		10'b1101000100: color_data = 12'b000000000000;
		10'b1101000101: color_data = 12'b000000000000;
		10'b1101000110: color_data = 12'b000000000000;
		10'b1101000111: color_data = 12'b000000000000;
		10'b1101001000: color_data = 12'b000000000000;
		10'b1101100011: color_data = 12'b000000000000;
		10'b1101100100: color_data = 12'b000000000000;
		10'b1101100101: color_data = 12'b000000000000;
		10'b1101100110: color_data = 12'b000000000000;
		10'b1101100111: color_data = 12'b000000000000;
		10'b1110000100: color_data = 12'b000000000000;
		10'b1110000101: color_data = 12'b000000000000;
		10'b1110000110: color_data = 12'b000000000000;
        default: color_data = 12'b111111111111;
	endcase
endmodule