module LRBack_rom (
	input wire clk,
    input wire [5:0] row,
    input wire [8:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 384 + col) >= 0 && (row * 384 + col) <= 420) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 439 && (row * 384 + col) <= 499) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 518 && (row * 384 + col) <= 801) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 827 && (row * 384 + col) <= 879) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 905 && (row * 384 + col) <= 1182) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 1191 && (row * 384 + col) <= 1204) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 1214 && (row * 384 + col) <= 1260) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 1270 && (row * 384 + col) <= 1283) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 1292 && (row * 384 + col) <= 1564) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 1571 && (row * 384 + col) <= 1594) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 1600 && (row * 384 + col) <= 1642) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 1648 && (row * 384 + col) <= 1671) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 1678 && (row * 384 + col) <= 1946) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 1952 && (row * 384 + col) <= 1980) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 1986 && (row * 384 + col) <= 2024) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 2030 && (row * 384 + col) <= 2058) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 2064 && (row * 384 + col) <= 2328) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 2334 && (row * 384 + col) <= 2366) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 2372 && (row * 384 + col) <= 2406) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 2412 && (row * 384 + col) <= 2444) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 2450 && (row * 384 + col) <= 2711) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 2716 && (row * 384 + col) <= 2752) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 2758 && (row * 384 + col) <= 2788) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 2794 && (row * 384 + col) <= 2830) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 2835 && (row * 384 + col) <= 3094) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 3099 && (row * 384 + col) <= 3101) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3102 && (row * 384 + col) <= 3104) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 3105 && (row * 384 + col) <= 3138) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3143 && (row * 384 + col) <= 3171) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 3176 && (row * 384 + col) <= 3201) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3202 && (row * 384 + col) <= 3210) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 3211 && (row * 384 + col) <= 3215) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3220 && (row * 384 + col) <= 3476) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 3481 && (row * 384 + col) <= 3485) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3486 && (row * 384 + col) <= 3488) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 3489 && (row * 384 + col) <= 3524) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3528 && (row * 384 + col) <= 3554) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 3558 && (row * 384 + col) <= 3585) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3586 && (row * 384 + col) <= 3594) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 3595 && (row * 384 + col) <= 3601) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3606 && (row * 384 + col) <= 3859) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 3864 && (row * 384 + col) <= 3869) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3870 && (row * 384 + col) <= 3872) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 3873 && (row * 384 + col) <= 3909) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3913 && (row * 384 + col) <= 3937) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 3941 && (row * 384 + col) <= 3969) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3970 && (row * 384 + col) <= 3978) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 3979 && (row * 384 + col) <= 3986) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 3991 && (row * 384 + col) <= 4242) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 4246 && (row * 384 + col) <= 4253) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4254 && (row * 384 + col) <= 4256) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 4257 && (row * 384 + col) <= 4294) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4298 && (row * 384 + col) <= 4320) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 4324 && (row * 384 + col) <= 4353) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4354 && (row * 384 + col) <= 4356) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 4357 && (row * 384 + col) <= 4362) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4363 && (row * 384 + col) <= 4365) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 4366 && (row * 384 + col) <= 4372) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4376 && (row * 384 + col) <= 4625) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 4629 && (row * 384 + col) <= 4637) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4638 && (row * 384 + col) <= 4640) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 4641 && (row * 384 + col) <= 4679) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4683 && (row * 384 + col) <= 4703) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 4707 && (row * 384 + col) <= 4737) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4738 && (row * 384 + col) <= 4740) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 4741 && (row * 384 + col) <= 4746) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4747 && (row * 384 + col) <= 4749) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 4750 && (row * 384 + col) <= 4757) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 4761 && (row * 384 + col) <= 5008) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5012 && (row * 384 + col) <= 5021) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5022 && (row * 384 + col) <= 5024) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 5025 && (row * 384 + col) <= 5061) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5067 && (row * 384 + col) <= 5087) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5093 && (row * 384 + col) <= 5121) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5122 && (row * 384 + col) <= 5124) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 5125 && (row * 384 + col) <= 5130) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5131 && (row * 384 + col) <= 5133) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 5134 && (row * 384 + col) <= 5142) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5146 && (row * 384 + col) <= 5391) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5395 && (row * 384 + col) <= 5405) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5406 && (row * 384 + col) <= 5408) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 5409 && (row * 384 + col) <= 5442) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5450 && (row * 384 + col) <= 5472) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5480 && (row * 384 + col) <= 5505) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5506 && (row * 384 + col) <= 5514) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 5515 && (row * 384 + col) <= 5527) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5531 && (row * 384 + col) <= 5774) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5778 && (row * 384 + col) <= 5789) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5790 && (row * 384 + col) <= 5792) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 5793 && (row * 384 + col) <= 5824) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5831 && (row * 384 + col) <= 5859) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5866 && (row * 384 + col) <= 5889) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5890 && (row * 384 + col) <= 5898) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 5899 && (row * 384 + col) <= 5912) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 5916 && (row * 384 + col) <= 5933) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5938 && (row * 384 + col) <= 5946) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5957 && (row * 384 + col) <= 5966) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5973 && (row * 384 + col) <= 5982) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 5990 && (row * 384 + col) <= 5996) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6000 && (row * 384 + col) <= 6006) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6010 && (row * 384 + col) <= 6020) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6036 && (row * 384 + col) <= 6040) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6048 && (row * 384 + col) <= 6065) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6076 && (row * 384 + col) <= 6079) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6095 && (row * 384 + col) <= 6099) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6106 && (row * 384 + col) <= 6112) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6123 && (row * 384 + col) <= 6127) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6143 && (row * 384 + col) <= 6157) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6161 && (row * 384 + col) <= 6173) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6174 && (row * 384 + col) <= 6176) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 6177 && (row * 384 + col) <= 6205) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6212 && (row * 384 + col) <= 6246) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6253 && (row * 384 + col) <= 6273) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6274 && (row * 384 + col) <= 6282) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 6283 && (row * 384 + col) <= 6297) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6301 && (row * 384 + col) <= 6317) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6322 && (row * 384 + col) <= 6330) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6341 && (row * 384 + col) <= 6350) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6357 && (row * 384 + col) <= 6366) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6374 && (row * 384 + col) <= 6380) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6384 && (row * 384 + col) <= 6390) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6394 && (row * 384 + col) <= 6404) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6420 && (row * 384 + col) <= 6424) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6432 && (row * 384 + col) <= 6449) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6460 && (row * 384 + col) <= 6463) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6479 && (row * 384 + col) <= 6483) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6490 && (row * 384 + col) <= 6496) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6507 && (row * 384 + col) <= 6511) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6527 && (row * 384 + col) <= 6540) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6544 && (row * 384 + col) <= 6557) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6558 && (row * 384 + col) <= 6560) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 6561 && (row * 384 + col) <= 6587) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6594 && (row * 384 + col) <= 6632) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6639 && (row * 384 + col) <= 6657) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6658 && (row * 384 + col) <= 6660) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 6661 && (row * 384 + col) <= 6663) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6664 && (row * 384 + col) <= 6666) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 6667 && (row * 384 + col) <= 6682) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6686 && (row * 384 + col) <= 6701) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6706 && (row * 384 + col) <= 6714) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6725 && (row * 384 + col) <= 6734) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6741 && (row * 384 + col) <= 6750) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6758 && (row * 384 + col) <= 6764) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6768 && (row * 384 + col) <= 6774) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6778 && (row * 384 + col) <= 6788) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6804 && (row * 384 + col) <= 6808) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6816 && (row * 384 + col) <= 6833) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6844 && (row * 384 + col) <= 6847) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6863 && (row * 384 + col) <= 6867) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6874 && (row * 384 + col) <= 6880) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6891 && (row * 384 + col) <= 6895) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6911 && (row * 384 + col) <= 6923) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 6927 && (row * 384 + col) <= 6941) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6942 && (row * 384 + col) <= 6944) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 6945 && (row * 384 + col) <= 6968) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 6975 && (row * 384 + col) <= 7019) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7026 && (row * 384 + col) <= 7041) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7042 && (row * 384 + col) <= 7044) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7045 && (row * 384 + col) <= 7047) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7048 && (row * 384 + col) <= 7050) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7051 && (row * 384 + col) <= 7067) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7071 && (row * 384 + col) <= 7085) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7090 && (row * 384 + col) <= 7098) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7102 && (row * 384 + col) <= 7108) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7112 && (row * 384 + col) <= 7115) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7119 && (row * 384 + col) <= 7124) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7128 && (row * 384 + col) <= 7131) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7135 && (row * 384 + col) <= 7141) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7145 && (row * 384 + col) <= 7148) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7152 && (row * 384 + col) <= 7154) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7159 && (row * 384 + col) <= 7178) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7182 && (row * 384 + col) <= 7189) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7193 && (row * 384 + col) <= 7199) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7203 && (row * 384 + col) <= 7214) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7218 && (row * 384 + col) <= 7237) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7241 && (row * 384 + col) <= 7248) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7252 && (row * 384 + col) <= 7257) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7261 && (row * 384 + col) <= 7264) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7268 && (row * 384 + col) <= 7274) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7278 && (row * 384 + col) <= 7285) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7289 && (row * 384 + col) <= 7306) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7310 && (row * 384 + col) <= 7325) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7326 && (row * 384 + col) <= 7328) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7329 && (row * 384 + col) <= 7349) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7357 && (row * 384 + col) <= 7405) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7413 && (row * 384 + col) <= 7425) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7426 && (row * 384 + col) <= 7428) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7429 && (row * 384 + col) <= 7431) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7432 && (row * 384 + col) <= 7434) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7435 && (row * 384 + col) <= 7452) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7456 && (row * 384 + col) <= 7482) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7486 && (row * 384 + col) <= 7492) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7496 && (row * 384 + col) <= 7499) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7503 && (row * 384 + col) <= 7508) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7512 && (row * 384 + col) <= 7515) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7519 && (row * 384 + col) <= 7525) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7529 && (row * 384 + col) <= 7532) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7536 && (row * 384 + col) <= 7538) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7543 && (row * 384 + col) <= 7562) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7566 && (row * 384 + col) <= 7573) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7577 && (row * 384 + col) <= 7583) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7587 && (row * 384 + col) <= 7598) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7602 && (row * 384 + col) <= 7621) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7625 && (row * 384 + col) <= 7632) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7636 && (row * 384 + col) <= 7641) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7645 && (row * 384 + col) <= 7648) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7652 && (row * 384 + col) <= 7658) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7662 && (row * 384 + col) <= 7669) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7673 && (row * 384 + col) <= 7689) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7693 && (row * 384 + col) <= 7709) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7710 && (row * 384 + col) <= 7721) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7722 && (row * 384 + col) <= 7730) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7738 && (row * 384 + col) <= 7792) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7800 && (row * 384 + col) <= 7809) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7810 && (row * 384 + col) <= 7812) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7813 && (row * 384 + col) <= 7818) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7819 && (row * 384 + col) <= 7821) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 7822 && (row * 384 + col) <= 7837) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 7841 && (row * 384 + col) <= 7866) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7870 && (row * 384 + col) <= 7876) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7880 && (row * 384 + col) <= 7883) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7887 && (row * 384 + col) <= 7892) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7896 && (row * 384 + col) <= 7899) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7903 && (row * 384 + col) <= 7909) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7913 && (row * 384 + col) <= 7916) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7920 && (row * 384 + col) <= 7922) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7927 && (row * 384 + col) <= 7946) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7950 && (row * 384 + col) <= 7957) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7961 && (row * 384 + col) <= 7967) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7971 && (row * 384 + col) <= 7982) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 7986 && (row * 384 + col) <= 8005) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8009 && (row * 384 + col) <= 8016) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8020 && (row * 384 + col) <= 8025) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8029 && (row * 384 + col) <= 8032) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8036 && (row * 384 + col) <= 8042) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8046 && (row * 384 + col) <= 8053) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8057 && (row * 384 + col) <= 8072) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8076 && (row * 384 + col) <= 8093) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8094 && (row * 384 + col) <= 8105) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 8106 && (row * 384 + col) <= 8111) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8119 && (row * 384 + col) <= 8147) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8151 && (row * 384 + col) <= 8179) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8187 && (row * 384 + col) <= 8193) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8194 && (row * 384 + col) <= 8196) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 8197 && (row * 384 + col) <= 8202) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8203 && (row * 384 + col) <= 8205) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 8206 && (row * 384 + col) <= 8222) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8226 && (row * 384 + col) <= 8250) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8254 && (row * 384 + col) <= 8260) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8264 && (row * 384 + col) <= 8267) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8271 && (row * 384 + col) <= 8276) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8280 && (row * 384 + col) <= 8283) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8287 && (row * 384 + col) <= 8293) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8297 && (row * 384 + col) <= 8300) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8304 && (row * 384 + col) <= 8306) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8311 && (row * 384 + col) <= 8330) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8334 && (row * 384 + col) <= 8341) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8345 && (row * 384 + col) <= 8351) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8355 && (row * 384 + col) <= 8366) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8370 && (row * 384 + col) <= 8389) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8393 && (row * 384 + col) <= 8400) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8404 && (row * 384 + col) <= 8409) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8413 && (row * 384 + col) <= 8416) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8420 && (row * 384 + col) <= 8426) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8430 && (row * 384 + col) <= 8437) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8441 && (row * 384 + col) <= 8456) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8459 && (row * 384 + col) <= 8477) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8478 && (row * 384 + col) <= 8489) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 8490 && (row * 384 + col) <= 8493) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8500 && (row * 384 + col) <= 8531) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8535 && (row * 384 + col) <= 8566) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8573 && (row * 384 + col) <= 8577) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8578 && (row * 384 + col) <= 8580) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 8581 && (row * 384 + col) <= 8586) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8587 && (row * 384 + col) <= 8589) color_data <= 12'b101010101010; else
        if ((row * 384 + col) >= 8590 && (row * 384 + col) <= 8607) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8610 && (row * 384 + col) <= 8634) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8645 && (row * 384 + col) <= 8651) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8664 && (row * 384 + col) <= 8667) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8671 && (row * 384 + col) <= 8684) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8691 && (row * 384 + col) <= 8714) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8718 && (row * 384 + col) <= 8725) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8729 && (row * 384 + col) <= 8735) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8739 && (row * 384 + col) <= 8753) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8761 && (row * 384 + col) <= 8773) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8777 && (row * 384 + col) <= 8784) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8797 && (row * 384 + col) <= 8800) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8811 && (row * 384 + col) <= 8821) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8825 && (row * 384 + col) <= 8839) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8843 && (row * 384 + col) <= 8874) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8881 && (row * 384 + col) <= 8915) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8919 && (row * 384 + col) <= 8953) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 8960 && (row * 384 + col) <= 8991) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 8995 && (row * 384 + col) <= 9018) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9029 && (row * 384 + col) <= 9035) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9048 && (row * 384 + col) <= 9051) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9055 && (row * 384 + col) <= 9068) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9075 && (row * 384 + col) <= 9098) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9102 && (row * 384 + col) <= 9109) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9113 && (row * 384 + col) <= 9119) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9123 && (row * 384 + col) <= 9137) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9145 && (row * 384 + col) <= 9157) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9161 && (row * 384 + col) <= 9168) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9181 && (row * 384 + col) <= 9184) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9195 && (row * 384 + col) <= 9205) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9209 && (row * 384 + col) <= 9222) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9226 && (row * 384 + col) <= 9256) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 9263 && (row * 384 + col) <= 9299) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9303 && (row * 384 + col) <= 9339) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9346 && (row * 384 + col) <= 9376) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 9380 && (row * 384 + col) <= 9402) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9413 && (row * 384 + col) <= 9419) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9432 && (row * 384 + col) <= 9435) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9439 && (row * 384 + col) <= 9452) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9459 && (row * 384 + col) <= 9482) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9486 && (row * 384 + col) <= 9493) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9497 && (row * 384 + col) <= 9503) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9507 && (row * 384 + col) <= 9521) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9529 && (row * 384 + col) <= 9541) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9545 && (row * 384 + col) <= 9552) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9565 && (row * 384 + col) <= 9568) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9579 && (row * 384 + col) <= 9589) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9593 && (row * 384 + col) <= 9606) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9610 && (row * 384 + col) <= 9638) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 9644 && (row * 384 + col) <= 9683) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9687 && (row * 384 + col) <= 9726) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9732 && (row * 384 + col) <= 9760) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 9764 && (row * 384 + col) <= 9786) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9790 && (row * 384 + col) <= 9796) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9800 && (row * 384 + col) <= 9803) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9807 && (row * 384 + col) <= 9812) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9816 && (row * 384 + col) <= 9819) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9823 && (row * 384 + col) <= 9829) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9833 && (row * 384 + col) <= 9836) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9840 && (row * 384 + col) <= 9842) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9847 && (row * 384 + col) <= 9866) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9870 && (row * 384 + col) <= 9877) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9881 && (row * 384 + col) <= 9887) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9891 && (row * 384 + col) <= 9912) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9916 && (row * 384 + col) <= 9925) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9929 && (row * 384 + col) <= 9936) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9940 && (row * 384 + col) <= 9945) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9949 && (row * 384 + col) <= 9952) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9956 && (row * 384 + col) <= 9959) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9963 && (row * 384 + col) <= 9973) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9977 && (row * 384 + col) <= 9989) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 9993 && (row * 384 + col) <= 10020) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 10026 && (row * 384 + col) <= 10067) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10071 && (row * 384 + col) <= 10112) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10118 && (row * 384 + col) <= 10145) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 10149 && (row * 384 + col) <= 10170) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10174 && (row * 384 + col) <= 10180) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10184 && (row * 384 + col) <= 10187) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10191 && (row * 384 + col) <= 10196) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10200 && (row * 384 + col) <= 10203) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10207 && (row * 384 + col) <= 10213) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10217 && (row * 384 + col) <= 10220) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10224 && (row * 384 + col) <= 10226) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10231 && (row * 384 + col) <= 10250) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10254 && (row * 384 + col) <= 10261) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10265 && (row * 384 + col) <= 10271) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10275 && (row * 384 + col) <= 10296) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10300 && (row * 384 + col) <= 10309) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10313 && (row * 384 + col) <= 10320) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10324 && (row * 384 + col) <= 10329) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10333 && (row * 384 + col) <= 10336) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10340 && (row * 384 + col) <= 10343) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10347 && (row * 384 + col) <= 10357) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10361 && (row * 384 + col) <= 10373) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10376 && (row * 384 + col) <= 10401) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 10408 && (row * 384 + col) <= 10444) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10461 && (row * 384 + col) <= 10498) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10505 && (row * 384 + col) <= 10530) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 10533 && (row * 384 + col) <= 10541) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10546 && (row * 384 + col) <= 10554) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10558 && (row * 384 + col) <= 10564) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10568 && (row * 384 + col) <= 10571) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10575 && (row * 384 + col) <= 10580) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10584 && (row * 384 + col) <= 10587) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10591 && (row * 384 + col) <= 10597) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10601 && (row * 384 + col) <= 10604) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10608 && (row * 384 + col) <= 10610) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10615 && (row * 384 + col) <= 10634) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10638 && (row * 384 + col) <= 10645) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10649 && (row * 384 + col) <= 10655) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10659 && (row * 384 + col) <= 10680) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10684 && (row * 384 + col) <= 10693) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10697 && (row * 384 + col) <= 10704) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10708 && (row * 384 + col) <= 10713) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10717 && (row * 384 + col) <= 10720) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10724 && (row * 384 + col) <= 10727) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10731 && (row * 384 + col) <= 10741) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10745 && (row * 384 + col) <= 10757) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10760 && (row * 384 + col) <= 10783) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 10790 && (row * 384 + col) <= 10828) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10845 && (row * 384 + col) <= 10884) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10891 && (row * 384 + col) <= 10914) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 10917 && (row * 384 + col) <= 10925) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10930 && (row * 384 + col) <= 10938) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10949 && (row * 384 + col) <= 10955) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10959 && (row * 384 + col) <= 10964) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10968 && (row * 384 + col) <= 10974) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10982 && (row * 384 + col) <= 10988) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 10992 && (row * 384 + col) <= 10998) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11002 && (row * 384 + col) <= 11018) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11022 && (row * 384 + col) <= 11032) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11040 && (row * 384 + col) <= 11054) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11065 && (row * 384 + col) <= 11077) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11081 && (row * 384 + col) <= 11088) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11092 && (row * 384 + col) <= 11097) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11101 && (row * 384 + col) <= 11104) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11108 && (row * 384 + col) <= 11114) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11118 && (row * 384 + col) <= 11125) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11129 && (row * 384 + col) <= 11140) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11144 && (row * 384 + col) <= 11164) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 11171 && (row * 384 + col) <= 11212) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11229 && (row * 384 + col) <= 11271) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11278 && (row * 384 + col) <= 11298) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 11302 && (row * 384 + col) <= 11309) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11314 && (row * 384 + col) <= 11322) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11333 && (row * 384 + col) <= 11339) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11343 && (row * 384 + col) <= 11348) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11352 && (row * 384 + col) <= 11358) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11366 && (row * 384 + col) <= 11372) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11376 && (row * 384 + col) <= 11382) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11386 && (row * 384 + col) <= 11402) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11406 && (row * 384 + col) <= 11416) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11424 && (row * 384 + col) <= 11438) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11449 && (row * 384 + col) <= 11461) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11465 && (row * 384 + col) <= 11472) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11476 && (row * 384 + col) <= 11481) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11485 && (row * 384 + col) <= 11488) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11492 && (row * 384 + col) <= 11498) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11502 && (row * 384 + col) <= 11509) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11513 && (row * 384 + col) <= 11524) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11527 && (row * 384 + col) <= 11546) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 11553 && (row * 384 + col) <= 11603) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11607 && (row * 384 + col) <= 11657) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11664 && (row * 384 + col) <= 11683) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 11686 && (row * 384 + col) <= 11693) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11698 && (row * 384 + col) <= 11706) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11717 && (row * 384 + col) <= 11723) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11727 && (row * 384 + col) <= 11732) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11736 && (row * 384 + col) <= 11742) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11750 && (row * 384 + col) <= 11756) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11760 && (row * 384 + col) <= 11766) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11770 && (row * 384 + col) <= 11786) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11790 && (row * 384 + col) <= 11800) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11808 && (row * 384 + col) <= 11822) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11833 && (row * 384 + col) <= 11845) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11849 && (row * 384 + col) <= 11856) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11860 && (row * 384 + col) <= 11865) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11869 && (row * 384 + col) <= 11872) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11876 && (row * 384 + col) <= 11882) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11886 && (row * 384 + col) <= 11893) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11897 && (row * 384 + col) <= 11907) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11911 && (row * 384 + col) <= 11928) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 11934 && (row * 384 + col) <= 11987) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 11991 && (row * 384 + col) <= 12044) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 12050 && (row * 384 + col) <= 12067) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 12071 && (row * 384 + col) <= 12291) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 12295 && (row * 384 + col) <= 12309) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 12316 && (row * 384 + col) <= 12371) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 12375 && (row * 384 + col) <= 12430) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 12437 && (row * 384 + col) <= 12451) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 12455 && (row * 384 + col) <= 12674) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 12678 && (row * 384 + col) <= 12691) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 12698 && (row * 384 + col) <= 12755) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 12759 && (row * 384 + col) <= 12816) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 12823 && (row * 384 + col) <= 12836) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 12840 && (row * 384 + col) <= 13058) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13062 && (row * 384 + col) <= 13073) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 13079 && (row * 384 + col) <= 13139) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13143 && (row * 384 + col) <= 13203) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13209 && (row * 384 + col) <= 13220) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 13224 && (row * 384 + col) <= 13442) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13445 && (row * 384 + col) <= 13455) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 13461 && (row * 384 + col) <= 13523) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13527 && (row * 384 + col) <= 13589) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13595 && (row * 384 + col) <= 13605) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 13608 && (row * 384 + col) <= 13825) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13829 && (row * 384 + col) <= 13837) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 13843 && (row * 384 + col) <= 13975) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 13981 && (row * 384 + col) <= 13989) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 13993 && (row * 384 + col) <= 14209) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 14212 && (row * 384 + col) <= 14219) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 14225 && (row * 384 + col) <= 14361) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 14367 && (row * 384 + col) <= 14374) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 14377 && (row * 384 + col) <= 14592) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 14596 && (row * 384 + col) <= 14601) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 14607 && (row * 384 + col) <= 14747) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 14753 && (row * 384 + col) <= 14758) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 14762 && (row * 384 + col) <= 14976) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 14980 && (row * 384 + col) <= 14983) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 14989 && (row * 384 + col) <= 15133) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 15139 && (row * 384 + col) <= 15142) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 15146 && (row * 384 + col) <= 15360) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 15363 && (row * 384 + col) <= 15366) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 15371 && (row * 384 + col) <= 15519) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 15524 && (row * 384 + col) <= 15527) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 15530 && (row * 384 + col) <= 15744) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 15747 && (row * 384 + col) <= 15748) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 15753 && (row * 384 + col) <= 15905) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 15910 && (row * 384 + col) <= 15911) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 15914 && (row * 384 + col) <= 16128) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 16131 && (row * 384 + col) <= 16131) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 16136 && (row * 384 + col) <= 16290) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 16295 && (row * 384 + col) <= 16295) color_data <= 12'b110011001100; else
        if ((row * 384 + col) >= 16298 && (row * 384 + col) <= 16512) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 16518 && (row * 384 + col) <= 16676) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 16682 && (row * 384 + col) <= 16897) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 16901 && (row * 384 + col) <= 17061) color_data <= 12'b111111111111; else
        if ((row * 384 + col) >= 17065 && (row * 384 + col) < 17664) color_data <= 12'b111111111111; else
        color_data <= 12'b000000000000;
    end
endmodule