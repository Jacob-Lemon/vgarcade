`timescale 1ns / 1ps
module xfill_rom (
    input wire clk,
    input wire [7:0] row,
    input wire [9:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 584 + col) >= 0 && (row * 584 + col) <= 40271) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 40272 && (row * 584 + col) <= 40275) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 40276 && (row * 584 + col) <= 40840) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 40841 && (row * 584 + col) <= 40861) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 40862 && (row * 584 + col) <= 41423) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 41424 && (row * 584 + col) <= 41446) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 41447 && (row * 584 + col) <= 42006) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 42007 && (row * 584 + col) <= 42031) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 42032 && (row * 584 + col) <= 42590) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 42591 && (row * 584 + col) <= 42616) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 42617 && (row * 584 + col) <= 43174) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 43175 && (row * 584 + col) <= 43201) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 43202 && (row * 584 + col) <= 43758) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 43759 && (row * 584 + col) <= 43785) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 43786 && (row * 584 + col) <= 44342) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 44343 && (row * 584 + col) <= 44370) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 44371 && (row * 584 + col) <= 44926) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 44927 && (row * 584 + col) <= 44954) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 44955 && (row * 584 + col) <= 45510) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 45511 && (row * 584 + col) <= 45539) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 45540 && (row * 584 + col) <= 46094) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 46095 && (row * 584 + col) <= 46123) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 46124 && (row * 584 + col) <= 46678) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 46679 && (row * 584 + col) <= 46707) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 46708 && (row * 584 + col) <= 47262) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 47263 && (row * 584 + col) <= 47292) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 47293 && (row * 584 + col) <= 47846) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 47847 && (row * 584 + col) <= 47876) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 47877 && (row * 584 + col) <= 48430) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 48431 && (row * 584 + col) <= 48460) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 48461 && (row * 584 + col) <= 49014) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 49015 && (row * 584 + col) <= 49044) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 49045 && (row * 584 + col) <= 49598) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 49599 && (row * 584 + col) <= 49629) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 49630 && (row * 584 + col) <= 50182) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 50183 && (row * 584 + col) <= 50213) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 50214 && (row * 584 + col) <= 50766) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 50767 && (row * 584 + col) <= 50797) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 50798 && (row * 584 + col) <= 51350) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 51351 && (row * 584 + col) <= 51381) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 51382 && (row * 584 + col) <= 51935) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 51936 && (row * 584 + col) <= 51966) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 51967 && (row * 584 + col) <= 52519) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 52520 && (row * 584 + col) <= 52550) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 52551 && (row * 584 + col) <= 53104) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 53105 && (row * 584 + col) <= 53134) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 53135 && (row * 584 + col) <= 53688) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 53689 && (row * 584 + col) <= 53718) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 53719 && (row * 584 + col) <= 54273) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 54274 && (row * 584 + col) <= 54302) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 54303 && (row * 584 + col) <= 54858) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 54859 && (row * 584 + col) <= 54886) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 54887 && (row * 584 + col) <= 55444) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 55445 && (row * 584 + col) <= 55470) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 55471 && (row * 584 + col) <= 56028) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 56029 && (row * 584 + col) <= 56054) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 56055 && (row * 584 + col) <= 56612) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 56613 && (row * 584 + col) <= 56639) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 56640 && (row * 584 + col) <= 57195) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 57196 && (row * 584 + col) <= 57223) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 57224 && (row * 584 + col) <= 57779) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 57780 && (row * 584 + col) <= 57807) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 57808 && (row * 584 + col) <= 58363) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 58364 && (row * 584 + col) <= 58391) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 58392 && (row * 584 + col) <= 58947) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 58948 && (row * 584 + col) <= 58975) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 58976 && (row * 584 + col) <= 59531) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 59532 && (row * 584 + col) <= 59559) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 59560 && (row * 584 + col) <= 60115) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 60116 && (row * 584 + col) <= 60143) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 60144 && (row * 584 + col) <= 60699) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 60700 && (row * 584 + col) <= 60727) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 60728 && (row * 584 + col) <= 61283) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 61284 && (row * 584 + col) <= 61311) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 61312 && (row * 584 + col) <= 61867) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 61868 && (row * 584 + col) <= 61895) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 61896 && (row * 584 + col) <= 62451) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 62452 && (row * 584 + col) <= 62479) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 62480 && (row * 584 + col) <= 63035) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 63036 && (row * 584 + col) <= 63063) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 63064 && (row * 584 + col) <= 63619) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 63620 && (row * 584 + col) <= 63647) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 63648 && (row * 584 + col) <= 64203) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 64204 && (row * 584 + col) <= 64231) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 64232 && (row * 584 + col) <= 64787) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 64788 && (row * 584 + col) <= 64815) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 64816 && (row * 584 + col) <= 65371) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 65372 && (row * 584 + col) <= 65399) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 65400 && (row * 584 + col) <= 65955) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 65956 && (row * 584 + col) <= 65983) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 65984 && (row * 584 + col) <= 66539) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 66540 && (row * 584 + col) <= 66567) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 66568 && (row * 584 + col) <= 67123) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 67124 && (row * 584 + col) <= 67151) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 67152 && (row * 584 + col) <= 67708) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 67709 && (row * 584 + col) <= 67735) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 67736 && (row * 584 + col) <= 68292) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 68293 && (row * 584 + col) <= 68318) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 68319 && (row * 584 + col) <= 68876) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 68877 && (row * 584 + col) <= 68902) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 68903 && (row * 584 + col) <= 69460) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 69461 && (row * 584 + col) <= 69486) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 69487 && (row * 584 + col) <= 70044) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 70045 && (row * 584 + col) <= 70070) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 70071 && (row * 584 + col) <= 70628) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 70629 && (row * 584 + col) <= 70654) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 70655 && (row * 584 + col) <= 71212) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 71213 && (row * 584 + col) <= 71238) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 71239 && (row * 584 + col) <= 71796) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 71797 && (row * 584 + col) <= 71822) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 71823 && (row * 584 + col) <= 72381) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 72382 && (row * 584 + col) <= 72406) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 72407 && (row * 584 + col) <= 72965) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 72966 && (row * 584 + col) <= 72989) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 72990 && (row * 584 + col) <= 73549) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 73550 && (row * 584 + col) <= 73573) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 73574 && (row * 584 + col) <= 74133) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 74134 && (row * 584 + col) <= 74157) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 74158 && (row * 584 + col) <= 74717) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 74718 && (row * 584 + col) <= 74741) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 74742 && (row * 584 + col) <= 75302) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 75303 && (row * 584 + col) <= 75324) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 75325 && (row * 584 + col) <= 75886) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 75887 && (row * 584 + col) <= 75908) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 75909 && (row * 584 + col) <= 76470) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 76471 && (row * 584 + col) <= 76492) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 76493 && (row * 584 + col) <= 77054) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 77055 && (row * 584 + col) <= 77076) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 77077 && (row * 584 + col) <= 77639) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 77640 && (row * 584 + col) <= 77659) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 77660 && (row * 584 + col) <= 78223) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 78224 && (row * 584 + col) <= 78243) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 78244 && (row * 584 + col) <= 78808) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 78809 && (row * 584 + col) <= 78827) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 78828 && (row * 584 + col) <= 79392) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 79393 && (row * 584 + col) <= 79410) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 79411 && (row * 584 + col) <= 79976) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 79977 && (row * 584 + col) <= 79994) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 79995 && (row * 584 + col) <= 80561) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 80562 && (row * 584 + col) <= 80577) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 80578 && (row * 584 + col) <= 81146) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 81147 && (row * 584 + col) <= 81161) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 81162 && (row * 584 + col) <= 81730) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 81731 && (row * 584 + col) <= 81744) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 81745 && (row * 584 + col) <= 82315) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 82316 && (row * 584 + col) <= 82327) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 82328 && (row * 584 + col) <= 82900) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 82901 && (row * 584 + col) <= 82910) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 82911 && (row * 584 + col) <= 83485) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 83486 && (row * 584 + col) <= 83493) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 83494 && (row * 584 + col) <= 84071) color_data <= 12'b000000000000; else
        if ((row * 584 + col) >= 84072 && (row * 584 + col) <= 84075) color_data <= 12'b111111111111; else
        if ((row * 584 + col) >= 84076 && (row * 584 + col) < 97528) color_data <= 12'b000000000000; else
        color_data <= 12'b000000000000;
    end
endmodule
