module player_shielded_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [6:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "distributed" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		14'b00000010100000: color_data = 12'b000000000000;
		14'b00000010100001: color_data = 12'b000000000000;
		14'b00000010100010: color_data = 12'b000000000000;
		14'b00000010100011: color_data = 12'b000000000000;
		14'b00000010100100: color_data = 12'b000000000000;
		14'b00000010100101: color_data = 12'b000000000000;
		14'b00000100011101: color_data = 12'b000000000000;
		14'b00000100011110: color_data = 12'b000000000000;
		14'b00000100011111: color_data = 12'b000000000000;
		14'b00000100100000: color_data = 12'b111111111010;
		14'b00000100100001: color_data = 12'b111111111010;
		14'b00000100100010: color_data = 12'b111111111010;
		14'b00000100100011: color_data = 12'b111111111010;
		14'b00000100100100: color_data = 12'b111111111010;
		14'b00000100100101: color_data = 12'b111111111010;
		14'b00000100100110: color_data = 12'b000000000000;
		14'b00000100100111: color_data = 12'b000000000000;
		14'b00000100101000: color_data = 12'b000000000000;
		14'b00000110011100: color_data = 12'b000000000000;
		14'b00000110011101: color_data = 12'b111111111010;
		14'b00000110011110: color_data = 12'b111111111010;
		14'b00000110011111: color_data = 12'b111111111010;
		14'b00000110100000: color_data = 12'b111111111010;
		14'b00000110100001: color_data = 12'b111111111010;
		14'b00000110100010: color_data = 12'b111111111010;
		14'b00000110100011: color_data = 12'b111111111010;
		14'b00000110100100: color_data = 12'b111111111010;
		14'b00000110100101: color_data = 12'b111111111010;
		14'b00000110100110: color_data = 12'b111111111010;
		14'b00000110100111: color_data = 12'b111111111010;
		14'b00000110101000: color_data = 12'b111111111010;
		14'b00000110101001: color_data = 12'b000000000000;
		14'b00001000011010: color_data = 12'b000000000000;
		14'b00001000011011: color_data = 12'b000000000000;
		14'b00001000011100: color_data = 12'b111111111010;
		14'b00001000011101: color_data = 12'b111111111010;
		14'b00001000011110: color_data = 12'b111111111010;
		14'b00001000011111: color_data = 12'b111111111010;
		14'b00001000100000: color_data = 12'b111111111010;
		14'b00001000100001: color_data = 12'b111111111010;
		14'b00001000100010: color_data = 12'b111111111010;
		14'b00001000100011: color_data = 12'b111111111010;
		14'b00001000100100: color_data = 12'b111111111010;
		14'b00001000100101: color_data = 12'b111111111010;
		14'b00001000100110: color_data = 12'b111111111010;
		14'b00001000100111: color_data = 12'b111111111010;
		14'b00001000101000: color_data = 12'b111111111010;
		14'b00001000101001: color_data = 12'b111111111010;
		14'b00001000101010: color_data = 12'b000000000000;
		14'b00001000101011: color_data = 12'b000000000000;
		14'b00001010011001: color_data = 12'b000000000000;
		14'b00001010011010: color_data = 12'b111111111010;
		14'b00001010011011: color_data = 12'b111111111010;
		14'b00001010011100: color_data = 12'b111111111010;
		14'b00001010011101: color_data = 12'b111111111010;
		14'b00001010011110: color_data = 12'b111111111010;
		14'b00001010011111: color_data = 12'b111111111010;
		14'b00001010100000: color_data = 12'b111111111010;
		14'b00001010100001: color_data = 12'b111111111010;
		14'b00001010100010: color_data = 12'b111111111010;
		14'b00001010100011: color_data = 12'b111111111010;
		14'b00001010100100: color_data = 12'b111111111010;
		14'b00001010100101: color_data = 12'b111111111010;
		14'b00001010100110: color_data = 12'b111111111010;
		14'b00001010100111: color_data = 12'b111111111010;
		14'b00001010101000: color_data = 12'b111111111010;
		14'b00001010101001: color_data = 12'b111111111010;
		14'b00001010101010: color_data = 12'b111111111010;
		14'b00001010101011: color_data = 12'b111111111010;
		14'b00001010101100: color_data = 12'b000000000000;
		14'b00001100011001: color_data = 12'b000000000000;
		14'b00001100011010: color_data = 12'b111111111010;
		14'b00001100011011: color_data = 12'b111111111010;
		14'b00001100011100: color_data = 12'b111111111010;
		14'b00001100011101: color_data = 12'b111111111010;
		14'b00001100011110: color_data = 12'b111111111010;
		14'b00001100011111: color_data = 12'b111111111010;
		14'b00001100100000: color_data = 12'b111111111010;
		14'b00001100100001: color_data = 12'b111111111010;
		14'b00001100100010: color_data = 12'b111111111010;
		14'b00001100100011: color_data = 12'b111111111010;
		14'b00001100100100: color_data = 12'b111111111010;
		14'b00001100100101: color_data = 12'b111111111010;
		14'b00001100100110: color_data = 12'b111111111010;
		14'b00001100100111: color_data = 12'b111111111010;
		14'b00001100101000: color_data = 12'b111111111010;
		14'b00001100101001: color_data = 12'b111111111010;
		14'b00001100101010: color_data = 12'b111111111010;
		14'b00001100101011: color_data = 12'b111111111010;
		14'b00001100101100: color_data = 12'b000000000000;
		14'b00001110011000: color_data = 12'b000000000000;
		14'b00001110011001: color_data = 12'b111111111010;
		14'b00001110011010: color_data = 12'b111111111010;
		14'b00001110011011: color_data = 12'b111111111010;
		14'b00001110011100: color_data = 12'b111111111010;
		14'b00001110011101: color_data = 12'b111111111010;
		14'b00001110011110: color_data = 12'b111111111010;
		14'b00001110011111: color_data = 12'b111111111010;
		14'b00001110100000: color_data = 12'b111111111010;
		14'b00001110100001: color_data = 12'b111111111010;
		14'b00001110100010: color_data = 12'b111111111010;
		14'b00001110100011: color_data = 12'b111111111010;
		14'b00001110100100: color_data = 12'b111111111010;
		14'b00001110100101: color_data = 12'b111111111010;
		14'b00001110100110: color_data = 12'b111111111010;
		14'b00001110100111: color_data = 12'b111111111010;
		14'b00001110101000: color_data = 12'b111111111010;
		14'b00001110101001: color_data = 12'b111111111010;
		14'b00001110101010: color_data = 12'b111111111010;
		14'b00001110101011: color_data = 12'b111111111010;
		14'b00001110101100: color_data = 12'b111111111010;
		14'b00001110101101: color_data = 12'b000000000000;
		14'b00001110101110: color_data = 12'b000000000000;
		14'b00010000011000: color_data = 12'b000000000000;
		14'b00010000011001: color_data = 12'b000000000000;
		14'b00010000011010: color_data = 12'b000000000000;
		14'b00010000011011: color_data = 12'b000000000000;
		14'b00010000011100: color_data = 12'b000000000000;
		14'b00010000011101: color_data = 12'b000000000000;
		14'b00010000011110: color_data = 12'b000000000000;
		14'b00010000011111: color_data = 12'b000000000000;
		14'b00010000100000: color_data = 12'b000000000000;
		14'b00010000100001: color_data = 12'b000000000000;
		14'b00010000100010: color_data = 12'b000000000000;
		14'b00010000100011: color_data = 12'b000000000000;
		14'b00010000100100: color_data = 12'b000000000000;
		14'b00010000100101: color_data = 12'b000000000000;
		14'b00010000100110: color_data = 12'b000000000000;
		14'b00010000100111: color_data = 12'b000000000000;
		14'b00010000101000: color_data = 12'b000000000000;
		14'b00010000101001: color_data = 12'b000000000000;
		14'b00010000101010: color_data = 12'b000000000000;
		14'b00010000101011: color_data = 12'b000000000000;
		14'b00010000101100: color_data = 12'b000000000000;
		14'b00010000101101: color_data = 12'b000000000000;
		14'b00010000101110: color_data = 12'b000000000000;
		14'b00010010010111: color_data = 12'b000000000000;
		14'b00010010011000: color_data = 12'b111111111010;
		14'b00010010011001: color_data = 12'b111111111010;
		14'b00010010011010: color_data = 12'b111111111010;
		14'b00010010011011: color_data = 12'b000000000000;
		14'b00010010011100: color_data = 12'b111011101110;
		14'b00010010011101: color_data = 12'b111011101110;
		14'b00010010011110: color_data = 12'b111011101110;
		14'b00010010011111: color_data = 12'b111011101110;
		14'b00010010100000: color_data = 12'b111011101110;
		14'b00010010100001: color_data = 12'b111011101110;
		14'b00010010100010: color_data = 12'b000000000000;
		14'b00010010100011: color_data = 12'b111111111010;
		14'b00010010100100: color_data = 12'b111111111010;
		14'b00010010100101: color_data = 12'b000000000000;
		14'b00010010100110: color_data = 12'b111011101110;
		14'b00010010100111: color_data = 12'b111011101110;
		14'b00010010101000: color_data = 12'b111011101110;
		14'b00010010101001: color_data = 12'b111011101110;
		14'b00010010101010: color_data = 12'b111011101110;
		14'b00010010101011: color_data = 12'b000000000000;
		14'b00010010101100: color_data = 12'b111111111010;
		14'b00010010101101: color_data = 12'b111111111010;
		14'b00010010101110: color_data = 12'b000000000000;
		14'b00010100010111: color_data = 12'b000000000000;
		14'b00010100011000: color_data = 12'b111111111010;
		14'b00010100011001: color_data = 12'b111111111010;
		14'b00010100011010: color_data = 12'b111111111010;
		14'b00010100011011: color_data = 12'b000000000000;
		14'b00010100011100: color_data = 12'b111011101110;
		14'b00010100011101: color_data = 12'b111011101110;
		14'b00010100011110: color_data = 12'b111011101110;
		14'b00010100011111: color_data = 12'b001101001100;
		14'b00010100100000: color_data = 12'b001101001100;
		14'b00010100100001: color_data = 12'b111011101110;
		14'b00010100100010: color_data = 12'b000000000000;
		14'b00010100100011: color_data = 12'b111111111010;
		14'b00010100100100: color_data = 12'b111111111010;
		14'b00010100100101: color_data = 12'b000000000000;
		14'b00010100100110: color_data = 12'b111011101110;
		14'b00010100100111: color_data = 12'b001101001100;
		14'b00010100101000: color_data = 12'b001101001100;
		14'b00010100101001: color_data = 12'b111011101110;
		14'b00010100101010: color_data = 12'b111011101110;
		14'b00010100101011: color_data = 12'b000000000000;
		14'b00010100101100: color_data = 12'b111111111010;
		14'b00010100101101: color_data = 12'b111111111010;
		14'b00010100101110: color_data = 12'b000000000000;
		14'b00010110010110: color_data = 12'b000000000000;
		14'b00010110010111: color_data = 12'b111111111010;
		14'b00010110011000: color_data = 12'b111111111010;
		14'b00010110011001: color_data = 12'b111111111010;
		14'b00010110011010: color_data = 12'b111111111010;
		14'b00010110011011: color_data = 12'b000000000000;
		14'b00010110011100: color_data = 12'b111011101110;
		14'b00010110011101: color_data = 12'b111011101110;
		14'b00010110011110: color_data = 12'b111011101110;
		14'b00010110011111: color_data = 12'b001101001100;
		14'b00010110100000: color_data = 12'b001101001100;
		14'b00010110100001: color_data = 12'b111011101110;
		14'b00010110100010: color_data = 12'b000000000000;
		14'b00010110100011: color_data = 12'b111111111010;
		14'b00010110100100: color_data = 12'b111111111010;
		14'b00010110100101: color_data = 12'b000000000000;
		14'b00010110100110: color_data = 12'b111011101110;
		14'b00010110100111: color_data = 12'b001101001100;
		14'b00010110101000: color_data = 12'b001101001100;
		14'b00010110101001: color_data = 12'b111011101110;
		14'b00010110101010: color_data = 12'b111011101110;
		14'b00010110101011: color_data = 12'b000000000000;
		14'b00010110101100: color_data = 12'b111111111010;
		14'b00010110101101: color_data = 12'b111111111010;
		14'b00010110101110: color_data = 12'b111111111010;
		14'b00010110101111: color_data = 12'b000000000000;
		14'b00011000010110: color_data = 12'b000000000000;
		14'b00011000010111: color_data = 12'b111111111010;
		14'b00011000011000: color_data = 12'b111111111010;
		14'b00011000011001: color_data = 12'b111111111010;
		14'b00011000011010: color_data = 12'b111111111010;
		14'b00011000011011: color_data = 12'b000000000000;
		14'b00011000011100: color_data = 12'b000000000000;
		14'b00011000011101: color_data = 12'b000000000000;
		14'b00011000011110: color_data = 12'b000000000000;
		14'b00011000011111: color_data = 12'b000000000000;
		14'b00011000100000: color_data = 12'b000000000000;
		14'b00011000100001: color_data = 12'b000000000000;
		14'b00011000100010: color_data = 12'b000000000000;
		14'b00011000100011: color_data = 12'b111111111010;
		14'b00011000100100: color_data = 12'b111111111010;
		14'b00011000100101: color_data = 12'b000000000000;
		14'b00011000100110: color_data = 12'b000000000000;
		14'b00011000100111: color_data = 12'b000000000000;
		14'b00011000101000: color_data = 12'b000000000000;
		14'b00011000101001: color_data = 12'b000000000000;
		14'b00011000101010: color_data = 12'b000000000000;
		14'b00011000101011: color_data = 12'b000000000000;
		14'b00011000101100: color_data = 12'b111111111010;
		14'b00011000101101: color_data = 12'b111111111010;
		14'b00011000101110: color_data = 12'b111111111010;
		14'b00011000101111: color_data = 12'b000000000000;
		14'b00011010010110: color_data = 12'b000000000000;
		14'b00011010010111: color_data = 12'b111111111010;
		14'b00011010011000: color_data = 12'b111111111010;
		14'b00011010011001: color_data = 12'b111111111010;
		14'b00011010011010: color_data = 12'b111111111010;
		14'b00011010011011: color_data = 12'b111111111010;
		14'b00011010011100: color_data = 12'b111111111010;
		14'b00011010011101: color_data = 12'b111111111010;
		14'b00011010011110: color_data = 12'b111111111010;
		14'b00011010011111: color_data = 12'b111111111010;
		14'b00011010100000: color_data = 12'b111111111010;
		14'b00011010100001: color_data = 12'b111111111010;
		14'b00011010100010: color_data = 12'b111111111010;
		14'b00011010100011: color_data = 12'b111111111010;
		14'b00011010100100: color_data = 12'b111111111010;
		14'b00011010100101: color_data = 12'b111111111010;
		14'b00011010100110: color_data = 12'b111111111010;
		14'b00011010100111: color_data = 12'b111111111010;
		14'b00011010101000: color_data = 12'b111111111010;
		14'b00011010101001: color_data = 12'b111111111010;
		14'b00011010101010: color_data = 12'b111111111010;
		14'b00011010101011: color_data = 12'b111111111010;
		14'b00011010101100: color_data = 12'b111111111010;
		14'b00011010101101: color_data = 12'b111111111010;
		14'b00011010101110: color_data = 12'b111111111010;
		14'b00011010101111: color_data = 12'b000000000000;
		14'b00011100010110: color_data = 12'b000000000000;
		14'b00011100010111: color_data = 12'b111111111010;
		14'b00011100011000: color_data = 12'b111111111010;
		14'b00011100011001: color_data = 12'b111111111010;
		14'b00011100011010: color_data = 12'b111111111010;
		14'b00011100011011: color_data = 12'b111111111010;
		14'b00011100011100: color_data = 12'b111111111010;
		14'b00011100011101: color_data = 12'b111111111010;
		14'b00011100011110: color_data = 12'b111111111010;
		14'b00011100011111: color_data = 12'b111111111010;
		14'b00011100100000: color_data = 12'b111111111010;
		14'b00011100100001: color_data = 12'b111111111010;
		14'b00011100100010: color_data = 12'b111111111010;
		14'b00011100100011: color_data = 12'b111111111010;
		14'b00011100100100: color_data = 12'b111111111010;
		14'b00011100100101: color_data = 12'b111111111010;
		14'b00011100100110: color_data = 12'b111111111010;
		14'b00011100100111: color_data = 12'b111111111010;
		14'b00011100101000: color_data = 12'b111111111010;
		14'b00011100101001: color_data = 12'b111111111010;
		14'b00011100101010: color_data = 12'b111111111010;
		14'b00011100101011: color_data = 12'b111111111010;
		14'b00011100101100: color_data = 12'b111111111010;
		14'b00011100101101: color_data = 12'b111111111010;
		14'b00011100101110: color_data = 12'b111111111010;
		14'b00011100101111: color_data = 12'b000000000000;
		14'b00011110010110: color_data = 12'b000000000000;
		14'b00011110010111: color_data = 12'b111111111010;
		14'b00011110011000: color_data = 12'b111111111010;
		14'b00011110011001: color_data = 12'b111111111010;
		14'b00011110011010: color_data = 12'b111111111010;
		14'b00011110011011: color_data = 12'b111111111010;
		14'b00011110011100: color_data = 12'b111111111010;
		14'b00011110011101: color_data = 12'b111111111010;
		14'b00011110011110: color_data = 12'b111111111010;
		14'b00011110011111: color_data = 12'b111111111010;
		14'b00011110100000: color_data = 12'b111111111010;
		14'b00011110100001: color_data = 12'b111111111010;
		14'b00011110100010: color_data = 12'b111111111010;
		14'b00011110100011: color_data = 12'b111111111010;
		14'b00011110100100: color_data = 12'b111111111010;
		14'b00011110100101: color_data = 12'b111111111010;
		14'b00011110100110: color_data = 12'b111111111010;
		14'b00011110100111: color_data = 12'b111111111010;
		14'b00011110101000: color_data = 12'b111111111010;
		14'b00011110101001: color_data = 12'b111111111010;
		14'b00011110101010: color_data = 12'b111111111010;
		14'b00011110101011: color_data = 12'b111111111010;
		14'b00011110101100: color_data = 12'b111111111010;
		14'b00011110101101: color_data = 12'b111111111010;
		14'b00011110101110: color_data = 12'b111111111010;
		14'b00011110101111: color_data = 12'b000000000000;
		14'b00100000010110: color_data = 12'b000000000000;
		14'b00100000010111: color_data = 12'b111111111010;
		14'b00100000011000: color_data = 12'b111111111010;
		14'b00100000011001: color_data = 12'b111111111010;
		14'b00100000011010: color_data = 12'b111111111010;
		14'b00100000011011: color_data = 12'b111111111010;
		14'b00100000011100: color_data = 12'b111111111010;
		14'b00100000011101: color_data = 12'b111111111010;
		14'b00100000011110: color_data = 12'b111111111010;
		14'b00100000011111: color_data = 12'b111111111010;
		14'b00100000100000: color_data = 12'b111111111010;
		14'b00100000100001: color_data = 12'b111111111010;
		14'b00100000100010: color_data = 12'b111111111010;
		14'b00100000100011: color_data = 12'b111111111010;
		14'b00100000100100: color_data = 12'b111111111010;
		14'b00100000100101: color_data = 12'b111111111010;
		14'b00100000100110: color_data = 12'b111111111010;
		14'b00100000100111: color_data = 12'b111111111010;
		14'b00100000101000: color_data = 12'b111111111010;
		14'b00100000101001: color_data = 12'b111111111010;
		14'b00100000101010: color_data = 12'b111111111010;
		14'b00100000101011: color_data = 12'b111111111010;
		14'b00100000101100: color_data = 12'b111111111010;
		14'b00100000101101: color_data = 12'b111111111010;
		14'b00100000101110: color_data = 12'b111111111010;
		14'b00100000101111: color_data = 12'b000000000000;
		14'b00100000111010: color_data = 12'b011101110111;
		14'b00100010010111: color_data = 12'b000000000000;
		14'b00100010011000: color_data = 12'b111111111010;
		14'b00100010011001: color_data = 12'b111111111010;
		14'b00100010011010: color_data = 12'b111111111010;
		14'b00100010011011: color_data = 12'b111111111010;
		14'b00100010011100: color_data = 12'b111111111010;
		14'b00100010011101: color_data = 12'b111111111010;
		14'b00100010011110: color_data = 12'b111111111010;
		14'b00100010011111: color_data = 12'b111111111010;
		14'b00100010100000: color_data = 12'b111111111010;
		14'b00100010100001: color_data = 12'b111111111010;
		14'b00100010100010: color_data = 12'b111111111010;
		14'b00100010100011: color_data = 12'b111111111010;
		14'b00100010100100: color_data = 12'b111111111010;
		14'b00100010100101: color_data = 12'b111111111010;
		14'b00100010100110: color_data = 12'b111111111010;
		14'b00100010100111: color_data = 12'b111111111010;
		14'b00100010101000: color_data = 12'b111111111010;
		14'b00100010101001: color_data = 12'b111111111010;
		14'b00100010101010: color_data = 12'b111111111010;
		14'b00100010101011: color_data = 12'b111111111010;
		14'b00100010101100: color_data = 12'b111111111010;
		14'b00100010101101: color_data = 12'b111111111010;
		14'b00100010101110: color_data = 12'b000000000000;
		14'b00100010111000: color_data = 12'b011101110111;
		14'b00100010111001: color_data = 12'b011101110111;
		14'b00100010111010: color_data = 12'b110011001100;
		14'b00100010111011: color_data = 12'b011101110111;
		14'b00100010111100: color_data = 12'b011101110111;
		14'b00100100010111: color_data = 12'b000000000000;
		14'b00100100011000: color_data = 12'b111111111010;
		14'b00100100011001: color_data = 12'b111111111010;
		14'b00100100011010: color_data = 12'b111111111010;
		14'b00100100011011: color_data = 12'b111111111010;
		14'b00100100011100: color_data = 12'b000000000000;
		14'b00100100011101: color_data = 12'b000000000000;
		14'b00100100011110: color_data = 12'b000000000000;
		14'b00100100011111: color_data = 12'b000000000000;
		14'b00100100100000: color_data = 12'b000000000000;
		14'b00100100100001: color_data = 12'b000000000000;
		14'b00100100100010: color_data = 12'b000000000000;
		14'b00100100100011: color_data = 12'b000000000000;
		14'b00100100100100: color_data = 12'b000000000000;
		14'b00100100100101: color_data = 12'b000000000000;
		14'b00100100100110: color_data = 12'b000000000000;
		14'b00100100100111: color_data = 12'b000000000000;
		14'b00100100101000: color_data = 12'b111111111010;
		14'b00100100101001: color_data = 12'b111111111010;
		14'b00100100101010: color_data = 12'b111111111010;
		14'b00100100101011: color_data = 12'b111111111010;
		14'b00100100101100: color_data = 12'b111111111010;
		14'b00100100101101: color_data = 12'b111111111010;
		14'b00100100101110: color_data = 12'b000000000000;
		14'b00100100110110: color_data = 12'b011101110111;
		14'b00100100110111: color_data = 12'b011101110111;
		14'b00100100111000: color_data = 12'b110011001100;
		14'b00100100111001: color_data = 12'b110011001100;
		14'b00100100111010: color_data = 12'b110011001100;
		14'b00100100111011: color_data = 12'b110011001100;
		14'b00100100111100: color_data = 12'b110011001100;
		14'b00100100111101: color_data = 12'b011101110111;
		14'b00100100111110: color_data = 12'b011101110111;
		14'b00100110010111: color_data = 12'b000000000000;
		14'b00100110011000: color_data = 12'b111111111010;
		14'b00100110011001: color_data = 12'b111111111010;
		14'b00100110011010: color_data = 12'b111111111010;
		14'b00100110011011: color_data = 12'b111111111010;
		14'b00100110011100: color_data = 12'b000000000000;
		14'b00100110011101: color_data = 12'b000000000000;
		14'b00100110011110: color_data = 12'b111011101110;
		14'b00100110011111: color_data = 12'b111011101110;
		14'b00100110100000: color_data = 12'b111011101110;
		14'b00100110100001: color_data = 12'b111011101110;
		14'b00100110100010: color_data = 12'b111011101110;
		14'b00100110100011: color_data = 12'b111011101110;
		14'b00100110100100: color_data = 12'b111011101110;
		14'b00100110100101: color_data = 12'b111011101110;
		14'b00100110100110: color_data = 12'b000000000000;
		14'b00100110100111: color_data = 12'b000000000000;
		14'b00100110101000: color_data = 12'b111111111010;
		14'b00100110101001: color_data = 12'b111111111010;
		14'b00100110101010: color_data = 12'b111111111010;
		14'b00100110101011: color_data = 12'b111111111010;
		14'b00100110101100: color_data = 12'b111111111010;
		14'b00100110101101: color_data = 12'b111111111010;
		14'b00100110101110: color_data = 12'b000000000000;
		14'b00100110110101: color_data = 12'b011101110111;
		14'b00100110110110: color_data = 12'b110011001100;
		14'b00100110110111: color_data = 12'b110011001100;
		14'b00100110111000: color_data = 12'b110011001100;
		14'b00100110111001: color_data = 12'b110011001100;
		14'b00100110111010: color_data = 12'b110011001100;
		14'b00100110111011: color_data = 12'b110011001100;
		14'b00100110111100: color_data = 12'b110011001100;
		14'b00100110111101: color_data = 12'b110011001100;
		14'b00100110111110: color_data = 12'b110011001100;
		14'b00100110111111: color_data = 12'b011101110111;
		14'b00101000011000: color_data = 12'b000000000000;
		14'b00101000011001: color_data = 12'b111111111010;
		14'b00101000011010: color_data = 12'b111111111010;
		14'b00101000011011: color_data = 12'b111111111010;
		14'b00101000011100: color_data = 12'b111111111010;
		14'b00101000011101: color_data = 12'b000000000000;
		14'b00101000011110: color_data = 12'b000000000000;
		14'b00101000011111: color_data = 12'b111011101110;
		14'b00101000100000: color_data = 12'b111011101110;
		14'b00101000100001: color_data = 12'b111011101110;
		14'b00101000100010: color_data = 12'b111011101110;
		14'b00101000100011: color_data = 12'b111011101110;
		14'b00101000100100: color_data = 12'b111011101110;
		14'b00101000100101: color_data = 12'b111011101110;
		14'b00101000100110: color_data = 12'b000000000000;
		14'b00101000100111: color_data = 12'b111111111010;
		14'b00101000101000: color_data = 12'b111111111010;
		14'b00101000101001: color_data = 12'b111111111010;
		14'b00101000101010: color_data = 12'b111111111010;
		14'b00101000101011: color_data = 12'b111111111010;
		14'b00101000101100: color_data = 12'b111111111010;
		14'b00101000101101: color_data = 12'b000000000000;
		14'b00101000110011: color_data = 12'b011101110111;
		14'b00101000110100: color_data = 12'b011101110111;
		14'b00101000110101: color_data = 12'b110011001100;
		14'b00101000110110: color_data = 12'b110011001100;
		14'b00101000110111: color_data = 12'b110011001100;
		14'b00101000111000: color_data = 12'b110011001100;
		14'b00101000111001: color_data = 12'b110011001100;
		14'b00101000111010: color_data = 12'b011101110111;
		14'b00101000111011: color_data = 12'b110011001100;
		14'b00101000111100: color_data = 12'b110011001100;
		14'b00101000111101: color_data = 12'b110011001100;
		14'b00101000111110: color_data = 12'b110011001100;
		14'b00101000111111: color_data = 12'b110011001100;
		14'b00101001000000: color_data = 12'b011101110111;
		14'b00101001000001: color_data = 12'b011101110111;
		14'b00101010011001: color_data = 12'b000000000000;
		14'b00101010011010: color_data = 12'b111111111010;
		14'b00101010011011: color_data = 12'b111111111010;
		14'b00101010011100: color_data = 12'b111111111010;
		14'b00101010011101: color_data = 12'b111111111010;
		14'b00101010011110: color_data = 12'b000000000000;
		14'b00101010011111: color_data = 12'b000000000000;
		14'b00101010100000: color_data = 12'b000000000000;
		14'b00101010100001: color_data = 12'b000000000000;
		14'b00101010100010: color_data = 12'b111011101110;
		14'b00101010100011: color_data = 12'b111011101110;
		14'b00101010100100: color_data = 12'b111011101110;
		14'b00101010100101: color_data = 12'b000000000000;
		14'b00101010100110: color_data = 12'b000000000000;
		14'b00101010100111: color_data = 12'b111111111010;
		14'b00101010101000: color_data = 12'b111111111010;
		14'b00101010101001: color_data = 12'b111111111010;
		14'b00101010101010: color_data = 12'b111111111010;
		14'b00101010101011: color_data = 12'b111111111010;
		14'b00101010101100: color_data = 12'b000000000000;
		14'b00101010110001: color_data = 12'b011101110111;
		14'b00101010110010: color_data = 12'b011101110111;
		14'b00101010110011: color_data = 12'b110011001100;
		14'b00101010110100: color_data = 12'b110011001100;
		14'b00101010110101: color_data = 12'b110011001100;
		14'b00101010110110: color_data = 12'b110011001100;
		14'b00101010110111: color_data = 12'b110011001100;
		14'b00101010111000: color_data = 12'b110011001100;
		14'b00101010111001: color_data = 12'b110011001100;
		14'b00101010111010: color_data = 12'b110011001100;
		14'b00101010111011: color_data = 12'b110011001100;
		14'b00101010111100: color_data = 12'b110011001100;
		14'b00101010111101: color_data = 12'b110011001100;
		14'b00101010111110: color_data = 12'b110011001100;
		14'b00101010111111: color_data = 12'b110011001100;
		14'b00101011000000: color_data = 12'b110011001100;
		14'b00101011000001: color_data = 12'b110011001100;
		14'b00101011000010: color_data = 12'b011101110111;
		14'b00101011000011: color_data = 12'b011101110111;
		14'b00101100011001: color_data = 12'b000000000000;
		14'b00101100011010: color_data = 12'b111111111010;
		14'b00101100011011: color_data = 12'b111111111010;
		14'b00101100011100: color_data = 12'b111111111010;
		14'b00101100011101: color_data = 12'b111111111010;
		14'b00101100011110: color_data = 12'b111111111010;
		14'b00101100011111: color_data = 12'b111111111010;
		14'b00101100100000: color_data = 12'b111111111010;
		14'b00101100100001: color_data = 12'b000000000000;
		14'b00101100100010: color_data = 12'b000000000000;
		14'b00101100100011: color_data = 12'b000000000000;
		14'b00101100100100: color_data = 12'b000000000000;
		14'b00101100100101: color_data = 12'b000000000000;
		14'b00101100100110: color_data = 12'b111111111010;
		14'b00101100100111: color_data = 12'b111111111010;
		14'b00101100101000: color_data = 12'b111111111010;
		14'b00101100101001: color_data = 12'b111111111010;
		14'b00101100101010: color_data = 12'b111111111010;
		14'b00101100101011: color_data = 12'b111111111010;
		14'b00101100101100: color_data = 12'b000000000000;
		14'b00101100101111: color_data = 12'b011101110111;
		14'b00101100110000: color_data = 12'b011101110111;
		14'b00101100110001: color_data = 12'b110011001100;
		14'b00101100110010: color_data = 12'b110011001100;
		14'b00101100110011: color_data = 12'b110011001100;
		14'b00101100110100: color_data = 12'b110011001100;
		14'b00101100110101: color_data = 12'b110011001100;
		14'b00101100110110: color_data = 12'b110011001100;
		14'b00101100110111: color_data = 12'b110011001100;
		14'b00101100111000: color_data = 12'b110011001100;
		14'b00101100111001: color_data = 12'b110011001100;
		14'b00101100111010: color_data = 12'b110011001100;
		14'b00101100111011: color_data = 12'b110011001100;
		14'b00101100111100: color_data = 12'b110011001100;
		14'b00101100111101: color_data = 12'b110011001100;
		14'b00101100111110: color_data = 12'b110011001100;
		14'b00101100111111: color_data = 12'b110011001100;
		14'b00101101000000: color_data = 12'b110011001100;
		14'b00101101000001: color_data = 12'b110011001100;
		14'b00101101000010: color_data = 12'b110011001100;
		14'b00101101000011: color_data = 12'b110011001100;
		14'b00101101000100: color_data = 12'b011101110111;
		14'b00101101000101: color_data = 12'b011101110111;
		14'b00101110011010: color_data = 12'b000000000000;
		14'b00101110011011: color_data = 12'b000000000000;
		14'b00101110011100: color_data = 12'b111111111010;
		14'b00101110011101: color_data = 12'b111111111010;
		14'b00101110011110: color_data = 12'b111111111010;
		14'b00101110011111: color_data = 12'b111111111010;
		14'b00101110100000: color_data = 12'b111111111010;
		14'b00101110100001: color_data = 12'b111111111010;
		14'b00101110100010: color_data = 12'b111111111010;
		14'b00101110100011: color_data = 12'b111111111010;
		14'b00101110100100: color_data = 12'b111111111010;
		14'b00101110100101: color_data = 12'b111111111010;
		14'b00101110100110: color_data = 12'b111111111010;
		14'b00101110100111: color_data = 12'b111111111010;
		14'b00101110101000: color_data = 12'b111111111010;
		14'b00101110101001: color_data = 12'b111111111010;
		14'b00101110101010: color_data = 12'b000000000000;
		14'b00101110101011: color_data = 12'b000000000000;
		14'b00101110101110: color_data = 12'b011101110111;
		14'b00101110101111: color_data = 12'b110011001100;
		14'b00101110110000: color_data = 12'b110011001100;
		14'b00101110110001: color_data = 12'b110011001100;
		14'b00101110110010: color_data = 12'b110011001100;
		14'b00101110110011: color_data = 12'b110011001100;
		14'b00101110110100: color_data = 12'b110011001100;
		14'b00101110110101: color_data = 12'b110011001100;
		14'b00101110110110: color_data = 12'b110011001100;
		14'b00101110110111: color_data = 12'b110011001100;
		14'b00101110111000: color_data = 12'b110011001100;
		14'b00101110111001: color_data = 12'b110011001100;
		14'b00101110111010: color_data = 12'b110011001100;
		14'b00101110111011: color_data = 12'b110011001100;
		14'b00101110111100: color_data = 12'b110011001100;
		14'b00101110111101: color_data = 12'b110011001100;
		14'b00101110111110: color_data = 12'b110011001100;
		14'b00101110111111: color_data = 12'b110011001100;
		14'b00101111000000: color_data = 12'b110011001100;
		14'b00101111000001: color_data = 12'b110011001100;
		14'b00101111000010: color_data = 12'b110011001100;
		14'b00101111000011: color_data = 12'b110011001100;
		14'b00101111000100: color_data = 12'b110011001100;
		14'b00101111000101: color_data = 12'b110011001100;
		14'b00101111000110: color_data = 12'b011101110111;
		14'b00110000011100: color_data = 12'b000000000000;
		14'b00110000011101: color_data = 12'b111111111010;
		14'b00110000011110: color_data = 12'b111111111010;
		14'b00110000011111: color_data = 12'b111111111010;
		14'b00110000100000: color_data = 12'b111111111010;
		14'b00110000100001: color_data = 12'b111111111010;
		14'b00110000100010: color_data = 12'b111111111010;
		14'b00110000100011: color_data = 12'b111111111010;
		14'b00110000100100: color_data = 12'b111111111010;
		14'b00110000100101: color_data = 12'b111111111010;
		14'b00110000100110: color_data = 12'b111111111010;
		14'b00110000100111: color_data = 12'b111111111010;
		14'b00110000101000: color_data = 12'b111111111010;
		14'b00110000101001: color_data = 12'b000000000000;
		14'b00110000101100: color_data = 12'b011101110111;
		14'b00110000101101: color_data = 12'b011101110111;
		14'b00110000101110: color_data = 12'b110011001100;
		14'b00110000101111: color_data = 12'b110011001100;
		14'b00110000110000: color_data = 12'b110011001100;
		14'b00110000110001: color_data = 12'b110011001100;
		14'b00110000110010: color_data = 12'b110011001100;
		14'b00110000110011: color_data = 12'b110011001100;
		14'b00110000110100: color_data = 12'b110011001100;
		14'b00110000110101: color_data = 12'b110011001100;
		14'b00110000110110: color_data = 12'b110011001100;
		14'b00110000110111: color_data = 12'b110011001100;
		14'b00110000111000: color_data = 12'b110011001100;
		14'b00110000111001: color_data = 12'b110011001100;
		14'b00110000111010: color_data = 12'b110011001100;
		14'b00110000111011: color_data = 12'b110011001100;
		14'b00110000111100: color_data = 12'b110011001100;
		14'b00110000111101: color_data = 12'b110011001100;
		14'b00110000111110: color_data = 12'b110011001100;
		14'b00110000111111: color_data = 12'b110011001100;
		14'b00110001000000: color_data = 12'b110011001100;
		14'b00110001000001: color_data = 12'b110011001100;
		14'b00110001000010: color_data = 12'b110011001100;
		14'b00110001000011: color_data = 12'b110011001100;
		14'b00110001000100: color_data = 12'b110011001100;
		14'b00110001000101: color_data = 12'b110011001100;
		14'b00110001000110: color_data = 12'b110011001100;
		14'b00110001000111: color_data = 12'b011101110111;
		14'b00110001001000: color_data = 12'b011101110111;
		14'b00110010011101: color_data = 12'b000000000000;
		14'b00110010011110: color_data = 12'b111111111010;
		14'b00110010011111: color_data = 12'b111111111010;
		14'b00110010100000: color_data = 12'b111111111010;
		14'b00110010100001: color_data = 12'b111111111010;
		14'b00110010100010: color_data = 12'b111111111010;
		14'b00110010100011: color_data = 12'b111111111010;
		14'b00110010100100: color_data = 12'b111111111010;
		14'b00110010100101: color_data = 12'b111111111010;
		14'b00110010100110: color_data = 12'b111111111010;
		14'b00110010100111: color_data = 12'b111111111010;
		14'b00110010101000: color_data = 12'b000000000000;
		14'b00110010101010: color_data = 12'b011101110111;
		14'b00110010101011: color_data = 12'b011101110111;
		14'b00110010101100: color_data = 12'b110011001100;
		14'b00110010101101: color_data = 12'b110011001100;
		14'b00110010101110: color_data = 12'b110011001100;
		14'b00110010101111: color_data = 12'b110011001100;
		14'b00110010110000: color_data = 12'b110011001100;
		14'b00110010110001: color_data = 12'b110011001100;
		14'b00110010110010: color_data = 12'b110011001100;
		14'b00110010110011: color_data = 12'b110011001100;
		14'b00110010110100: color_data = 12'b110011001100;
		14'b00110010110101: color_data = 12'b110011001100;
		14'b00110010110110: color_data = 12'b110011001100;
		14'b00110010110111: color_data = 12'b110011001100;
		14'b00110010111000: color_data = 12'b110011001100;
		14'b00110010111001: color_data = 12'b110011001100;
		14'b00110010111010: color_data = 12'b110011001100;
		14'b00110010111011: color_data = 12'b110011001100;
		14'b00110010111100: color_data = 12'b110011001100;
		14'b00110010111101: color_data = 12'b110011001100;
		14'b00110010111110: color_data = 12'b110011001100;
		14'b00110010111111: color_data = 12'b110011001100;
		14'b00110011000000: color_data = 12'b110011001100;
		14'b00110011000001: color_data = 12'b110011001100;
		14'b00110011000010: color_data = 12'b110011001100;
		14'b00110011000011: color_data = 12'b110011001100;
		14'b00110011000100: color_data = 12'b110011001100;
		14'b00110011000101: color_data = 12'b110011001100;
		14'b00110011000110: color_data = 12'b110011001100;
		14'b00110011000111: color_data = 12'b110011001100;
		14'b00110011001000: color_data = 12'b110011001100;
		14'b00110011001001: color_data = 12'b011101110111;
		14'b00110011001010: color_data = 12'b011101110111;
		14'b00110100000001: color_data = 12'b000000000000;
		14'b00110100000010: color_data = 12'b000000000000;
		14'b00110100000011: color_data = 12'b000000000000;
		14'b00110100000100: color_data = 12'b000000000000;
		14'b00110100000101: color_data = 12'b000000000000;
		14'b00110100000110: color_data = 12'b000000000000;
		14'b00110100000111: color_data = 12'b000000000000;
		14'b00110100001000: color_data = 12'b000000000000;
		14'b00110100001001: color_data = 12'b000000000000;
		14'b00110100001010: color_data = 12'b000000000000;
		14'b00110100001011: color_data = 12'b000000000000;
		14'b00110100001100: color_data = 12'b000000000000;
		14'b00110100001101: color_data = 12'b000000000000;
		14'b00110100001110: color_data = 12'b000000000000;
		14'b00110100001111: color_data = 12'b000000000000;
		14'b00110100010000: color_data = 12'b000000000000;
		14'b00110100010001: color_data = 12'b000000000000;
		14'b00110100010010: color_data = 12'b000000000000;
		14'b00110100010011: color_data = 12'b000000000000;
		14'b00110100010100: color_data = 12'b000000000000;
		14'b00110100010101: color_data = 12'b000000000000;
		14'b00110100010110: color_data = 12'b000000000000;
		14'b00110100010111: color_data = 12'b000000000000;
		14'b00110100011000: color_data = 12'b000000000000;
		14'b00110100011001: color_data = 12'b000000000000;
		14'b00110100011010: color_data = 12'b000000000000;
		14'b00110100011011: color_data = 12'b000000000000;
		14'b00110100011100: color_data = 12'b000000000000;
		14'b00110100011101: color_data = 12'b000000000000;
		14'b00110100011110: color_data = 12'b000000000000;
		14'b00110100011111: color_data = 12'b111111111010;
		14'b00110100100000: color_data = 12'b111111111010;
		14'b00110100100001: color_data = 12'b111111111010;
		14'b00110100100010: color_data = 12'b111111111010;
		14'b00110100100011: color_data = 12'b111111111010;
		14'b00110100100100: color_data = 12'b111111111010;
		14'b00110100100101: color_data = 12'b111111111010;
		14'b00110100100110: color_data = 12'b111111111010;
		14'b00110100100111: color_data = 12'b000000000000;
		14'b00110100101000: color_data = 12'b000000000000;
		14'b00110100101001: color_data = 12'b011101110111;
		14'b00110100101010: color_data = 12'b110011001100;
		14'b00110100101011: color_data = 12'b110011001100;
		14'b00110100101100: color_data = 12'b110011001100;
		14'b00110100101101: color_data = 12'b110011001100;
		14'b00110100101110: color_data = 12'b110011001100;
		14'b00110100101111: color_data = 12'b110011001100;
		14'b00110100110000: color_data = 12'b110011001100;
		14'b00110100110001: color_data = 12'b110011001100;
		14'b00110100110010: color_data = 12'b110011001100;
		14'b00110100110011: color_data = 12'b110011001100;
		14'b00110100110100: color_data = 12'b110011001100;
		14'b00110100110101: color_data = 12'b110011001100;
		14'b00110100110110: color_data = 12'b111011101110;
		14'b00110100110111: color_data = 12'b111011101110;
		14'b00110100111000: color_data = 12'b111011101110;
		14'b00110100111001: color_data = 12'b110011001100;
		14'b00110100111010: color_data = 12'b110011001100;
		14'b00110100111011: color_data = 12'b110011001100;
		14'b00110100111100: color_data = 12'b110011001100;
		14'b00110100111101: color_data = 12'b110011001100;
		14'b00110100111110: color_data = 12'b110011001100;
		14'b00110100111111: color_data = 12'b110011001100;
		14'b00110101000000: color_data = 12'b110011001100;
		14'b00110101000001: color_data = 12'b110011001100;
		14'b00110101000010: color_data = 12'b110011001100;
		14'b00110101000011: color_data = 12'b110011001100;
		14'b00110101000100: color_data = 12'b110011001100;
		14'b00110101000101: color_data = 12'b110011001100;
		14'b00110101000110: color_data = 12'b110011001100;
		14'b00110101000111: color_data = 12'b110011001100;
		14'b00110101001000: color_data = 12'b110011001100;
		14'b00110101001001: color_data = 12'b110011001100;
		14'b00110101001010: color_data = 12'b110011001100;
		14'b00110101001011: color_data = 12'b011101110111;
		14'b00110110000001: color_data = 12'b000000000000;
		14'b00110110000010: color_data = 12'b111111111010;
		14'b00110110000011: color_data = 12'b111111111010;
		14'b00110110000100: color_data = 12'b111111111010;
		14'b00110110000101: color_data = 12'b111111111010;
		14'b00110110000110: color_data = 12'b111111111010;
		14'b00110110000111: color_data = 12'b111111111010;
		14'b00110110001000: color_data = 12'b111111111010;
		14'b00110110001001: color_data = 12'b111111111010;
		14'b00110110001010: color_data = 12'b111111111010;
		14'b00110110001011: color_data = 12'b111111111010;
		14'b00110110001100: color_data = 12'b111111111010;
		14'b00110110001101: color_data = 12'b111111111010;
		14'b00110110001110: color_data = 12'b111111111010;
		14'b00110110001111: color_data = 12'b111111111010;
		14'b00110110010000: color_data = 12'b111111111010;
		14'b00110110010001: color_data = 12'b111111111010;
		14'b00110110010010: color_data = 12'b111000010010;
		14'b00110110010011: color_data = 12'b111000010010;
		14'b00110110010100: color_data = 12'b111000010010;
		14'b00110110010101: color_data = 12'b111000010010;
		14'b00110110010110: color_data = 12'b111000010010;
		14'b00110110010111: color_data = 12'b111000010010;
		14'b00110110011000: color_data = 12'b111000010010;
		14'b00110110011001: color_data = 12'b111000010010;
		14'b00110110011010: color_data = 12'b111000010010;
		14'b00110110011011: color_data = 12'b111000010010;
		14'b00110110011100: color_data = 12'b111000010010;
		14'b00110110011101: color_data = 12'b111000010010;
		14'b00110110011110: color_data = 12'b111000010010;
		14'b00110110011111: color_data = 12'b111000010010;
		14'b00110110100000: color_data = 12'b111000010010;
		14'b00110110100001: color_data = 12'b111000010010;
		14'b00110110100010: color_data = 12'b111000010010;
		14'b00110110100011: color_data = 12'b111000010010;
		14'b00110110100100: color_data = 12'b111000010010;
		14'b00110110100101: color_data = 12'b111000010010;
		14'b00110110100110: color_data = 12'b111000010010;
		14'b00110110100111: color_data = 12'b111000010010;
		14'b00110110101000: color_data = 12'b111000010010;
		14'b00110110101001: color_data = 12'b011101110111;
		14'b00110110101010: color_data = 12'b110011001100;
		14'b00110110101011: color_data = 12'b110011001100;
		14'b00110110101100: color_data = 12'b110011001100;
		14'b00110110101101: color_data = 12'b011101110111;
		14'b00110110101110: color_data = 12'b110011001100;
		14'b00110110101111: color_data = 12'b110011001100;
		14'b00110110110000: color_data = 12'b110011001100;
		14'b00110110110001: color_data = 12'b110011001100;
		14'b00110110110010: color_data = 12'b110011001100;
		14'b00110110110011: color_data = 12'b110011001100;
		14'b00110110110100: color_data = 12'b111011101110;
		14'b00110110110101: color_data = 12'b111011101110;
		14'b00110110110110: color_data = 12'b111011101110;
		14'b00110110110111: color_data = 12'b111011101110;
		14'b00110110111000: color_data = 12'b111011101110;
		14'b00110110111001: color_data = 12'b110011001100;
		14'b00110110111010: color_data = 12'b110011001100;
		14'b00110110111011: color_data = 12'b110011001100;
		14'b00110110111100: color_data = 12'b110011001100;
		14'b00110110111101: color_data = 12'b110011001100;
		14'b00110110111110: color_data = 12'b110011001100;
		14'b00110110111111: color_data = 12'b110011001100;
		14'b00110111000000: color_data = 12'b110011001100;
		14'b00110111000001: color_data = 12'b110011001100;
		14'b00110111000010: color_data = 12'b110011001100;
		14'b00110111000011: color_data = 12'b110011001100;
		14'b00110111000100: color_data = 12'b110011001100;
		14'b00110111000101: color_data = 12'b110011001100;
		14'b00110111000110: color_data = 12'b110011001100;
		14'b00110111000111: color_data = 12'b110011001100;
		14'b00110111001000: color_data = 12'b110011001100;
		14'b00110111001001: color_data = 12'b110011001100;
		14'b00110111001010: color_data = 12'b110011001100;
		14'b00110111001011: color_data = 12'b011101110111;
		14'b00111000000001: color_data = 12'b000000000000;
		14'b00111000000010: color_data = 12'b111111111010;
		14'b00111000000011: color_data = 12'b111111111010;
		14'b00111000000100: color_data = 12'b111111111010;
		14'b00111000000101: color_data = 12'b111111111010;
		14'b00111000000110: color_data = 12'b111111111010;
		14'b00111000000111: color_data = 12'b111111111010;
		14'b00111000001000: color_data = 12'b111111111010;
		14'b00111000001001: color_data = 12'b111111111010;
		14'b00111000001010: color_data = 12'b111111111010;
		14'b00111000001011: color_data = 12'b111111111010;
		14'b00111000001100: color_data = 12'b111111111010;
		14'b00111000001101: color_data = 12'b111111111010;
		14'b00111000001110: color_data = 12'b111111111010;
		14'b00111000001111: color_data = 12'b111111111010;
		14'b00111000010000: color_data = 12'b111111111010;
		14'b00111000010001: color_data = 12'b111111111010;
		14'b00111000010010: color_data = 12'b111000010010;
		14'b00111000010011: color_data = 12'b111000010010;
		14'b00111000010100: color_data = 12'b111000010010;
		14'b00111000010101: color_data = 12'b111000010010;
		14'b00111000010110: color_data = 12'b111000010010;
		14'b00111000010111: color_data = 12'b111000010010;
		14'b00111000011000: color_data = 12'b111000010010;
		14'b00111000011001: color_data = 12'b111000010010;
		14'b00111000011010: color_data = 12'b111000010010;
		14'b00111000011011: color_data = 12'b111000010010;
		14'b00111000011100: color_data = 12'b111000010010;
		14'b00111000011101: color_data = 12'b111000010010;
		14'b00111000011110: color_data = 12'b111000010010;
		14'b00111000011111: color_data = 12'b111000010010;
		14'b00111000100000: color_data = 12'b111000010010;
		14'b00111000100001: color_data = 12'b111000010010;
		14'b00111000100010: color_data = 12'b111000010010;
		14'b00111000100011: color_data = 12'b111000010010;
		14'b00111000100100: color_data = 12'b111000010010;
		14'b00111000100101: color_data = 12'b111000010010;
		14'b00111000100110: color_data = 12'b111000010010;
		14'b00111000100111: color_data = 12'b111000010010;
		14'b00111000101000: color_data = 12'b111000010010;
		14'b00111000101001: color_data = 12'b011101110111;
		14'b00111000101010: color_data = 12'b110011001100;
		14'b00111000101011: color_data = 12'b110011001100;
		14'b00111000101100: color_data = 12'b110011001100;
		14'b00111000101101: color_data = 12'b110011001100;
		14'b00111000101110: color_data = 12'b110011001100;
		14'b00111000101111: color_data = 12'b110011001100;
		14'b00111000110000: color_data = 12'b110011001100;
		14'b00111000110001: color_data = 12'b110011001100;
		14'b00111000110010: color_data = 12'b111011101110;
		14'b00111000110011: color_data = 12'b111011101110;
		14'b00111000110100: color_data = 12'b111011101110;
		14'b00111000110101: color_data = 12'b111011101110;
		14'b00111000110110: color_data = 12'b111011101110;
		14'b00111000110111: color_data = 12'b111011101110;
		14'b00111000111000: color_data = 12'b110011001100;
		14'b00111000111001: color_data = 12'b110011001100;
		14'b00111000111010: color_data = 12'b110011001100;
		14'b00111000111011: color_data = 12'b110011001100;
		14'b00111000111100: color_data = 12'b110011001100;
		14'b00111000111101: color_data = 12'b110011001100;
		14'b00111000111110: color_data = 12'b110011001100;
		14'b00111000111111: color_data = 12'b110011001100;
		14'b00111001000000: color_data = 12'b110011001100;
		14'b00111001000001: color_data = 12'b110011001100;
		14'b00111001000010: color_data = 12'b110011001100;
		14'b00111001000011: color_data = 12'b110011001100;
		14'b00111001000100: color_data = 12'b110011001100;
		14'b00111001000101: color_data = 12'b110011001100;
		14'b00111001000110: color_data = 12'b110011001100;
		14'b00111001000111: color_data = 12'b110011001100;
		14'b00111001001000: color_data = 12'b011101110111;
		14'b00111001001001: color_data = 12'b110011001100;
		14'b00111001001010: color_data = 12'b110011001100;
		14'b00111001001011: color_data = 12'b011101110111;
		14'b00111010000001: color_data = 12'b000000000000;
		14'b00111010000010: color_data = 12'b111111111010;
		14'b00111010000011: color_data = 12'b111111111010;
		14'b00111010000100: color_data = 12'b111111111010;
		14'b00111010000101: color_data = 12'b111111111010;
		14'b00111010000110: color_data = 12'b111111111010;
		14'b00111010000111: color_data = 12'b111111111010;
		14'b00111010001000: color_data = 12'b111111111010;
		14'b00111010001001: color_data = 12'b111111111010;
		14'b00111010001010: color_data = 12'b111111111010;
		14'b00111010001011: color_data = 12'b111111111010;
		14'b00111010001100: color_data = 12'b111111111010;
		14'b00111010001101: color_data = 12'b111111111010;
		14'b00111010001110: color_data = 12'b111111111010;
		14'b00111010001111: color_data = 12'b111111111010;
		14'b00111010010000: color_data = 12'b111111111010;
		14'b00111010010001: color_data = 12'b111111111010;
		14'b00111010010010: color_data = 12'b111000010010;
		14'b00111010010011: color_data = 12'b111000010010;
		14'b00111010010100: color_data = 12'b111000010010;
		14'b00111010010101: color_data = 12'b111000010010;
		14'b00111010010110: color_data = 12'b111000010010;
		14'b00111010010111: color_data = 12'b111000010010;
		14'b00111010011000: color_data = 12'b111000010010;
		14'b00111010011001: color_data = 12'b111000010010;
		14'b00111010011010: color_data = 12'b111000010010;
		14'b00111010011011: color_data = 12'b111000010010;
		14'b00111010011100: color_data = 12'b111000010010;
		14'b00111010011101: color_data = 12'b111000010010;
		14'b00111010011110: color_data = 12'b111000010010;
		14'b00111010011111: color_data = 12'b111000010010;
		14'b00111010100000: color_data = 12'b111000010010;
		14'b00111010100001: color_data = 12'b111000010010;
		14'b00111010100010: color_data = 12'b111000010010;
		14'b00111010100011: color_data = 12'b111000010010;
		14'b00111010100100: color_data = 12'b111000010010;
		14'b00111010100101: color_data = 12'b111000010010;
		14'b00111010100110: color_data = 12'b111000010010;
		14'b00111010100111: color_data = 12'b111000010010;
		14'b00111010101000: color_data = 12'b111000010010;
		14'b00111010101001: color_data = 12'b011101110111;
		14'b00111010101010: color_data = 12'b110011001100;
		14'b00111010101011: color_data = 12'b110011001100;
		14'b00111010101100: color_data = 12'b110011001100;
		14'b00111010101101: color_data = 12'b110011001100;
		14'b00111010101110: color_data = 12'b110011001100;
		14'b00111010101111: color_data = 12'b110011001100;
		14'b00111010110000: color_data = 12'b110011001100;
		14'b00111010110001: color_data = 12'b111011101110;
		14'b00111010110010: color_data = 12'b111011101110;
		14'b00111010110011: color_data = 12'b111011101110;
		14'b00111010110100: color_data = 12'b111011101110;
		14'b00111010110101: color_data = 12'b111011101110;
		14'b00111010110110: color_data = 12'b111011101110;
		14'b00111010110111: color_data = 12'b110011001100;
		14'b00111010111000: color_data = 12'b110011001100;
		14'b00111010111001: color_data = 12'b110011001100;
		14'b00111010111010: color_data = 12'b110011001100;
		14'b00111010111011: color_data = 12'b110011001100;
		14'b00111010111100: color_data = 12'b110011001100;
		14'b00111010111101: color_data = 12'b110011001100;
		14'b00111010111110: color_data = 12'b110011001100;
		14'b00111010111111: color_data = 12'b110011001100;
		14'b00111011000000: color_data = 12'b110011001100;
		14'b00111011000001: color_data = 12'b110011001100;
		14'b00111011000010: color_data = 12'b110011001100;
		14'b00111011000011: color_data = 12'b110011001100;
		14'b00111011000100: color_data = 12'b110011001100;
		14'b00111011000101: color_data = 12'b110011001100;
		14'b00111011000110: color_data = 12'b110011001100;
		14'b00111011000111: color_data = 12'b110011001100;
		14'b00111011001000: color_data = 12'b110011001100;
		14'b00111011001001: color_data = 12'b110011001100;
		14'b00111011001010: color_data = 12'b110011001100;
		14'b00111011001011: color_data = 12'b011101110111;
		14'b00111100000001: color_data = 12'b000000000000;
		14'b00111100000010: color_data = 12'b111111111010;
		14'b00111100000011: color_data = 12'b111111111010;
		14'b00111100000100: color_data = 12'b111111111010;
		14'b00111100000101: color_data = 12'b111111111010;
		14'b00111100000110: color_data = 12'b111111111010;
		14'b00111100000111: color_data = 12'b111111111010;
		14'b00111100001000: color_data = 12'b111111111010;
		14'b00111100001001: color_data = 12'b111111111010;
		14'b00111100001010: color_data = 12'b111111111010;
		14'b00111100001011: color_data = 12'b111111111010;
		14'b00111100001100: color_data = 12'b111111111010;
		14'b00111100001101: color_data = 12'b111111111010;
		14'b00111100001110: color_data = 12'b111111111010;
		14'b00111100001111: color_data = 12'b111111111010;
		14'b00111100010000: color_data = 12'b111111111010;
		14'b00111100010001: color_data = 12'b111111111010;
		14'b00111100010010: color_data = 12'b111000010010;
		14'b00111100010011: color_data = 12'b111000010010;
		14'b00111100010100: color_data = 12'b111000010010;
		14'b00111100010101: color_data = 12'b111000010010;
		14'b00111100010110: color_data = 12'b111000010010;
		14'b00111100010111: color_data = 12'b111000010010;
		14'b00111100011000: color_data = 12'b111000010010;
		14'b00111100011001: color_data = 12'b111000010010;
		14'b00111100011010: color_data = 12'b111000010010;
		14'b00111100011011: color_data = 12'b111000010010;
		14'b00111100011100: color_data = 12'b111000010010;
		14'b00111100011101: color_data = 12'b111000010010;
		14'b00111100011110: color_data = 12'b111000010010;
		14'b00111100011111: color_data = 12'b111000010010;
		14'b00111100100000: color_data = 12'b111000010010;
		14'b00111100100001: color_data = 12'b111000010010;
		14'b00111100100010: color_data = 12'b111000010010;
		14'b00111100100011: color_data = 12'b111000010010;
		14'b00111100100100: color_data = 12'b111000010010;
		14'b00111100100101: color_data = 12'b111000010010;
		14'b00111100100110: color_data = 12'b111000010010;
		14'b00111100100111: color_data = 12'b111000010010;
		14'b00111100101000: color_data = 12'b111000010010;
		14'b00111100101001: color_data = 12'b011101110111;
		14'b00111100101010: color_data = 12'b110011001100;
		14'b00111100101011: color_data = 12'b110011001100;
		14'b00111100101100: color_data = 12'b110011001100;
		14'b00111100101101: color_data = 12'b110011001100;
		14'b00111100101110: color_data = 12'b110011001100;
		14'b00111100101111: color_data = 12'b110011001100;
		14'b00111100110000: color_data = 12'b110011001100;
		14'b00111100110001: color_data = 12'b111011101110;
		14'b00111100110010: color_data = 12'b111011101110;
		14'b00111100110011: color_data = 12'b111011101110;
		14'b00111100110100: color_data = 12'b111011101110;
		14'b00111100110101: color_data = 12'b111011101110;
		14'b00111100110110: color_data = 12'b110011001100;
		14'b00111100110111: color_data = 12'b110011001100;
		14'b00111100111000: color_data = 12'b110011001100;
		14'b00111100111001: color_data = 12'b110011001100;
		14'b00111100111010: color_data = 12'b110011001100;
		14'b00111100111011: color_data = 12'b110011001100;
		14'b00111100111100: color_data = 12'b110011001100;
		14'b00111100111101: color_data = 12'b110011001100;
		14'b00111100111110: color_data = 12'b110011001100;
		14'b00111100111111: color_data = 12'b110011001100;
		14'b00111101000000: color_data = 12'b110011001100;
		14'b00111101000001: color_data = 12'b110011001100;
		14'b00111101000010: color_data = 12'b110011001100;
		14'b00111101000011: color_data = 12'b110011001100;
		14'b00111101000100: color_data = 12'b110011001100;
		14'b00111101000101: color_data = 12'b110011001100;
		14'b00111101000110: color_data = 12'b110011001100;
		14'b00111101000111: color_data = 12'b110011001100;
		14'b00111101001000: color_data = 12'b110011001100;
		14'b00111101001001: color_data = 12'b110011001100;
		14'b00111101001010: color_data = 12'b110011001100;
		14'b00111101001011: color_data = 12'b011101110111;
		14'b00111110000001: color_data = 12'b000000000000;
		14'b00111110000010: color_data = 12'b111111111010;
		14'b00111110000011: color_data = 12'b111111111010;
		14'b00111110000100: color_data = 12'b111111111010;
		14'b00111110000101: color_data = 12'b111111111010;
		14'b00111110000110: color_data = 12'b111111111010;
		14'b00111110000111: color_data = 12'b111111111010;
		14'b00111110001000: color_data = 12'b111111111010;
		14'b00111110001001: color_data = 12'b111111111010;
		14'b00111110001010: color_data = 12'b111111111010;
		14'b00111110001011: color_data = 12'b111111111010;
		14'b00111110001100: color_data = 12'b111111111010;
		14'b00111110001101: color_data = 12'b111111111010;
		14'b00111110001110: color_data = 12'b111111111010;
		14'b00111110001111: color_data = 12'b111111111010;
		14'b00111110010000: color_data = 12'b111111111010;
		14'b00111110010001: color_data = 12'b111111111010;
		14'b00111110010010: color_data = 12'b111000010010;
		14'b00111110010011: color_data = 12'b111000010010;
		14'b00111110010100: color_data = 12'b111000010010;
		14'b00111110010101: color_data = 12'b111000010010;
		14'b00111110010110: color_data = 12'b111000010010;
		14'b00111110010111: color_data = 12'b111000010010;
		14'b00111110011000: color_data = 12'b111000010010;
		14'b00111110011001: color_data = 12'b111000010010;
		14'b00111110011010: color_data = 12'b111000010010;
		14'b00111110011011: color_data = 12'b111000010010;
		14'b00111110011100: color_data = 12'b111000010010;
		14'b00111110011101: color_data = 12'b111000010010;
		14'b00111110011110: color_data = 12'b111000010010;
		14'b00111110011111: color_data = 12'b111000010010;
		14'b00111110100000: color_data = 12'b111000010010;
		14'b00111110100001: color_data = 12'b111000010010;
		14'b00111110100010: color_data = 12'b111000010010;
		14'b00111110100011: color_data = 12'b111000010010;
		14'b00111110100100: color_data = 12'b111000010010;
		14'b00111110100101: color_data = 12'b111000010010;
		14'b00111110100110: color_data = 12'b111000010010;
		14'b00111110100111: color_data = 12'b111000010010;
		14'b00111110101000: color_data = 12'b111000010010;
		14'b00111110101001: color_data = 12'b011101110111;
		14'b00111110101010: color_data = 12'b110011001100;
		14'b00111110101011: color_data = 12'b110011001100;
		14'b00111110101100: color_data = 12'b110011001100;
		14'b00111110101101: color_data = 12'b110011001100;
		14'b00111110101110: color_data = 12'b110011001100;
		14'b00111110101111: color_data = 12'b110011001100;
		14'b00111110110000: color_data = 12'b111011101110;
		14'b00111110110001: color_data = 12'b111011101110;
		14'b00111110110010: color_data = 12'b111011101110;
		14'b00111110110011: color_data = 12'b111011101110;
		14'b00111110110100: color_data = 12'b111011101110;
		14'b00111110110101: color_data = 12'b110011001100;
		14'b00111110110110: color_data = 12'b110011001100;
		14'b00111110110111: color_data = 12'b110011001100;
		14'b00111110111000: color_data = 12'b110011001100;
		14'b00111110111001: color_data = 12'b110011001100;
		14'b00111110111010: color_data = 12'b110011001100;
		14'b00111110111011: color_data = 12'b110011001100;
		14'b00111110111100: color_data = 12'b110011001100;
		14'b00111110111101: color_data = 12'b110011001100;
		14'b00111110111110: color_data = 12'b110011001100;
		14'b00111110111111: color_data = 12'b110011001100;
		14'b00111111000000: color_data = 12'b110011001100;
		14'b00111111000001: color_data = 12'b110011001100;
		14'b00111111000010: color_data = 12'b110011001100;
		14'b00111111000011: color_data = 12'b110011001100;
		14'b00111111000100: color_data = 12'b110011001100;
		14'b00111111000101: color_data = 12'b110011001100;
		14'b00111111000110: color_data = 12'b110011001100;
		14'b00111111000111: color_data = 12'b110011001100;
		14'b00111111001000: color_data = 12'b110011001100;
		14'b00111111001001: color_data = 12'b110011001100;
		14'b00111111001010: color_data = 12'b110011001100;
		14'b00111111001011: color_data = 12'b011101110111;
		14'b01000000000001: color_data = 12'b000000000000;
		14'b01000000000010: color_data = 12'b000000000000;
		14'b01000000000011: color_data = 12'b000000000000;
		14'b01000000000100: color_data = 12'b000000000000;
		14'b01000000000101: color_data = 12'b000000000000;
		14'b01000000000110: color_data = 12'b000000000000;
		14'b01000000000111: color_data = 12'b000000000000;
		14'b01000000001000: color_data = 12'b000000000000;
		14'b01000000001001: color_data = 12'b000000000000;
		14'b01000000001010: color_data = 12'b000000000000;
		14'b01000000001011: color_data = 12'b000000000000;
		14'b01000000001100: color_data = 12'b000000000000;
		14'b01000000001101: color_data = 12'b000000000000;
		14'b01000000001110: color_data = 12'b000000000000;
		14'b01000000001111: color_data = 12'b000000000000;
		14'b01000000010000: color_data = 12'b000000000000;
		14'b01000000010001: color_data = 12'b000000000000;
		14'b01000000010010: color_data = 12'b000000000000;
		14'b01000000010011: color_data = 12'b000000000000;
		14'b01000000010100: color_data = 12'b000000000000;
		14'b01000000010101: color_data = 12'b000000000000;
		14'b01000000010110: color_data = 12'b000000000000;
		14'b01000000010111: color_data = 12'b000000000000;
		14'b01000000011000: color_data = 12'b111000010010;
		14'b01000000011001: color_data = 12'b111000010010;
		14'b01000000011010: color_data = 12'b111000010010;
		14'b01000000011011: color_data = 12'b111000010010;
		14'b01000000011100: color_data = 12'b111000010010;
		14'b01000000011101: color_data = 12'b111000010010;
		14'b01000000011110: color_data = 12'b111000010010;
		14'b01000000011111: color_data = 12'b111000010010;
		14'b01000000100000: color_data = 12'b111000010010;
		14'b01000000100001: color_data = 12'b111000010010;
		14'b01000000100010: color_data = 12'b111000010010;
		14'b01000000100011: color_data = 12'b111000010010;
		14'b01000000100100: color_data = 12'b111000010010;
		14'b01000000100101: color_data = 12'b111000010010;
		14'b01000000100110: color_data = 12'b111000010010;
		14'b01000000100111: color_data = 12'b111000010010;
		14'b01000000101000: color_data = 12'b111000010010;
		14'b01000000101001: color_data = 12'b011101110111;
		14'b01000000101010: color_data = 12'b110011001100;
		14'b01000000101011: color_data = 12'b110011001100;
		14'b01000000101100: color_data = 12'b110011001100;
		14'b01000000101101: color_data = 12'b110011001100;
		14'b01000000101110: color_data = 12'b110011001100;
		14'b01000000101111: color_data = 12'b110011001100;
		14'b01000000110000: color_data = 12'b111011101110;
		14'b01000000110001: color_data = 12'b111011101110;
		14'b01000000110010: color_data = 12'b111011101110;
		14'b01000000110011: color_data = 12'b110011001100;
		14'b01000000110100: color_data = 12'b110011001100;
		14'b01000000110101: color_data = 12'b110011001100;
		14'b01000000110110: color_data = 12'b110011001100;
		14'b01000000110111: color_data = 12'b110011001100;
		14'b01000000111000: color_data = 12'b110011001100;
		14'b01000000111001: color_data = 12'b110011001100;
		14'b01000000111010: color_data = 12'b110011001100;
		14'b01000000111011: color_data = 12'b110011001100;
		14'b01000000111100: color_data = 12'b110011001100;
		14'b01000000111101: color_data = 12'b110011001100;
		14'b01000000111110: color_data = 12'b110011001100;
		14'b01000000111111: color_data = 12'b110011001100;
		14'b01000001000000: color_data = 12'b110011001100;
		14'b01000001000001: color_data = 12'b110011001100;
		14'b01000001000010: color_data = 12'b110011001100;
		14'b01000001000011: color_data = 12'b110011001100;
		14'b01000001000100: color_data = 12'b110011001100;
		14'b01000001000101: color_data = 12'b110011001100;
		14'b01000001000110: color_data = 12'b110011001100;
		14'b01000001000111: color_data = 12'b110011001100;
		14'b01000001001000: color_data = 12'b110011001100;
		14'b01000001001001: color_data = 12'b110011001100;
		14'b01000001001010: color_data = 12'b110011001100;
		14'b01000001001011: color_data = 12'b011101110111;
		14'b01000010010111: color_data = 12'b000000000000;
		14'b01000010011000: color_data = 12'b111000010010;
		14'b01000010011001: color_data = 12'b111000010010;
		14'b01000010011010: color_data = 12'b111000010010;
		14'b01000010011011: color_data = 12'b111000010010;
		14'b01000010011100: color_data = 12'b111000010010;
		14'b01000010011101: color_data = 12'b111000010010;
		14'b01000010011110: color_data = 12'b111000010010;
		14'b01000010011111: color_data = 12'b111000010010;
		14'b01000010100000: color_data = 12'b111000010010;
		14'b01000010100001: color_data = 12'b111000010010;
		14'b01000010100010: color_data = 12'b111000010010;
		14'b01000010100011: color_data = 12'b111000010010;
		14'b01000010100100: color_data = 12'b111000010010;
		14'b01000010100101: color_data = 12'b111000010010;
		14'b01000010100110: color_data = 12'b111000010010;
		14'b01000010100111: color_data = 12'b111000010010;
		14'b01000010101000: color_data = 12'b111000010010;
		14'b01000010101001: color_data = 12'b011101110111;
		14'b01000010101010: color_data = 12'b110011001100;
		14'b01000010101011: color_data = 12'b110011001100;
		14'b01000010101100: color_data = 12'b110011001100;
		14'b01000010101101: color_data = 12'b110011001100;
		14'b01000010101110: color_data = 12'b110011001100;
		14'b01000010101111: color_data = 12'b111011101110;
		14'b01000010110000: color_data = 12'b111011101110;
		14'b01000010110001: color_data = 12'b111011101110;
		14'b01000010110010: color_data = 12'b111011101110;
		14'b01000010110011: color_data = 12'b110011001100;
		14'b01000010110100: color_data = 12'b110011001100;
		14'b01000010110101: color_data = 12'b110011001100;
		14'b01000010110110: color_data = 12'b110011001100;
		14'b01000010110111: color_data = 12'b110011001100;
		14'b01000010111000: color_data = 12'b110011001100;
		14'b01000010111001: color_data = 12'b110011001100;
		14'b01000010111010: color_data = 12'b110011001100;
		14'b01000010111011: color_data = 12'b110011001100;
		14'b01000010111100: color_data = 12'b110011001100;
		14'b01000010111101: color_data = 12'b110011001100;
		14'b01000010111110: color_data = 12'b110011001100;
		14'b01000010111111: color_data = 12'b110011001100;
		14'b01000011000000: color_data = 12'b110011001100;
		14'b01000011000001: color_data = 12'b110011001100;
		14'b01000011000010: color_data = 12'b110011001100;
		14'b01000011000011: color_data = 12'b110011001100;
		14'b01000011000100: color_data = 12'b110011001100;
		14'b01000011000101: color_data = 12'b110011001100;
		14'b01000011000110: color_data = 12'b110011001100;
		14'b01000011000111: color_data = 12'b110011001100;
		14'b01000011001000: color_data = 12'b110011001100;
		14'b01000011001001: color_data = 12'b110011001100;
		14'b01000011001010: color_data = 12'b110011001100;
		14'b01000011001011: color_data = 12'b011101110111;
		14'b01000100010111: color_data = 12'b000000000000;
		14'b01000100011000: color_data = 12'b111000010010;
		14'b01000100011001: color_data = 12'b111000010010;
		14'b01000100011010: color_data = 12'b111000010010;
		14'b01000100011011: color_data = 12'b111000010010;
		14'b01000100011100: color_data = 12'b111000010010;
		14'b01000100011101: color_data = 12'b111000010010;
		14'b01000100011110: color_data = 12'b111000010010;
		14'b01000100011111: color_data = 12'b111000010010;
		14'b01000100100000: color_data = 12'b111000010010;
		14'b01000100100001: color_data = 12'b111000010010;
		14'b01000100100010: color_data = 12'b111000010010;
		14'b01000100100011: color_data = 12'b111000010010;
		14'b01000100100100: color_data = 12'b111000010010;
		14'b01000100100101: color_data = 12'b111000010010;
		14'b01000100100110: color_data = 12'b111000010010;
		14'b01000100100111: color_data = 12'b111000010010;
		14'b01000100101000: color_data = 12'b111000010010;
		14'b01000100101001: color_data = 12'b011101110111;
		14'b01000100101010: color_data = 12'b110011001100;
		14'b01000100101011: color_data = 12'b110011001100;
		14'b01000100101100: color_data = 12'b110011001100;
		14'b01000100101101: color_data = 12'b110011001100;
		14'b01000100101110: color_data = 12'b110011001100;
		14'b01000100101111: color_data = 12'b111011101110;
		14'b01000100110000: color_data = 12'b111011101110;
		14'b01000100110001: color_data = 12'b110011001100;
		14'b01000100110010: color_data = 12'b110011001100;
		14'b01000100110011: color_data = 12'b110011001100;
		14'b01000100110100: color_data = 12'b110011001100;
		14'b01000100110101: color_data = 12'b110011001100;
		14'b01000100110110: color_data = 12'b110011001100;
		14'b01000100110111: color_data = 12'b110011001100;
		14'b01000100111000: color_data = 12'b110011001100;
		14'b01000100111001: color_data = 12'b110011001100;
		14'b01000100111010: color_data = 12'b110011001100;
		14'b01000100111011: color_data = 12'b110011001100;
		14'b01000100111100: color_data = 12'b110011001100;
		14'b01000100111101: color_data = 12'b110011001100;
		14'b01000100111110: color_data = 12'b110011001100;
		14'b01000100111111: color_data = 12'b110011001100;
		14'b01000101000000: color_data = 12'b110011001100;
		14'b01000101000001: color_data = 12'b110011001100;
		14'b01000101000010: color_data = 12'b110011001100;
		14'b01000101000011: color_data = 12'b110011001100;
		14'b01000101000100: color_data = 12'b110011001100;
		14'b01000101000101: color_data = 12'b110011001100;
		14'b01000101000110: color_data = 12'b110011001100;
		14'b01000101000111: color_data = 12'b110011001100;
		14'b01000101001000: color_data = 12'b110011001100;
		14'b01000101001001: color_data = 12'b110011001100;
		14'b01000101001010: color_data = 12'b110011001100;
		14'b01000101001011: color_data = 12'b011101110111;
		14'b01000110010111: color_data = 12'b000000000000;
		14'b01000110011000: color_data = 12'b111000010010;
		14'b01000110011001: color_data = 12'b111000010010;
		14'b01000110011010: color_data = 12'b111000010010;
		14'b01000110011011: color_data = 12'b111000010010;
		14'b01000110011100: color_data = 12'b111000010010;
		14'b01000110011101: color_data = 12'b111000010010;
		14'b01000110011110: color_data = 12'b111000010010;
		14'b01000110011111: color_data = 12'b111000010010;
		14'b01000110100000: color_data = 12'b111000010010;
		14'b01000110100001: color_data = 12'b111000010010;
		14'b01000110100010: color_data = 12'b111000010010;
		14'b01000110100011: color_data = 12'b111000010010;
		14'b01000110100100: color_data = 12'b111000010010;
		14'b01000110100101: color_data = 12'b111000010010;
		14'b01000110100110: color_data = 12'b111000010010;
		14'b01000110100111: color_data = 12'b111000010010;
		14'b01000110101000: color_data = 12'b111000010010;
		14'b01000110101001: color_data = 12'b011101110111;
		14'b01000110101010: color_data = 12'b110011001100;
		14'b01000110101011: color_data = 12'b110011001100;
		14'b01000110101100: color_data = 12'b110011001100;
		14'b01000110101101: color_data = 12'b110011001100;
		14'b01000110101110: color_data = 12'b110011001100;
		14'b01000110101111: color_data = 12'b111011101110;
		14'b01000110110000: color_data = 12'b110011001100;
		14'b01000110110001: color_data = 12'b110011001100;
		14'b01000110110010: color_data = 12'b110011001100;
		14'b01000110110011: color_data = 12'b110011001100;
		14'b01000110110100: color_data = 12'b110011001100;
		14'b01000110110101: color_data = 12'b110011001100;
		14'b01000110110110: color_data = 12'b110011001100;
		14'b01000110110111: color_data = 12'b110011001100;
		14'b01000110111000: color_data = 12'b110011001100;
		14'b01000110111001: color_data = 12'b110011001100;
		14'b01000110111010: color_data = 12'b110011001100;
		14'b01000110111011: color_data = 12'b110011001100;
		14'b01000110111100: color_data = 12'b110011001100;
		14'b01000110111101: color_data = 12'b110011001100;
		14'b01000110111110: color_data = 12'b110011001100;
		14'b01000110111111: color_data = 12'b110011001100;
		14'b01000111000000: color_data = 12'b110011001100;
		14'b01000111000001: color_data = 12'b110011001100;
		14'b01000111000010: color_data = 12'b110011001100;
		14'b01000111000011: color_data = 12'b110011001100;
		14'b01000111000100: color_data = 12'b110011001100;
		14'b01000111000101: color_data = 12'b110011001100;
		14'b01000111000110: color_data = 12'b110011001100;
		14'b01000111000111: color_data = 12'b110011001100;
		14'b01000111001000: color_data = 12'b110011001100;
		14'b01000111001001: color_data = 12'b110011001100;
		14'b01000111001010: color_data = 12'b110011001100;
		14'b01000111001011: color_data = 12'b011101110111;
		14'b01001000010111: color_data = 12'b000000000000;
		14'b01001000011000: color_data = 12'b111000010010;
		14'b01001000011001: color_data = 12'b111000010010;
		14'b01001000011010: color_data = 12'b111000010010;
		14'b01001000011011: color_data = 12'b111000010010;
		14'b01001000011100: color_data = 12'b111000010010;
		14'b01001000011101: color_data = 12'b111000010010;
		14'b01001000011110: color_data = 12'b111000010010;
		14'b01001000011111: color_data = 12'b111000010010;
		14'b01001000100000: color_data = 12'b111000010010;
		14'b01001000100001: color_data = 12'b111000010010;
		14'b01001000100010: color_data = 12'b111000010010;
		14'b01001000100011: color_data = 12'b111000010010;
		14'b01001000100100: color_data = 12'b111000010010;
		14'b01001000100101: color_data = 12'b111000010010;
		14'b01001000100110: color_data = 12'b111000010010;
		14'b01001000100111: color_data = 12'b111000010010;
		14'b01001000101000: color_data = 12'b111000010010;
		14'b01001000101001: color_data = 12'b011101110111;
		14'b01001000101010: color_data = 12'b110011001100;
		14'b01001000101011: color_data = 12'b110011001100;
		14'b01001000101100: color_data = 12'b110011001100;
		14'b01001000101101: color_data = 12'b110011001100;
		14'b01001000101110: color_data = 12'b110011001100;
		14'b01001000101111: color_data = 12'b110011001100;
		14'b01001000110000: color_data = 12'b110011001100;
		14'b01001000110001: color_data = 12'b110011001100;
		14'b01001000110010: color_data = 12'b110011001100;
		14'b01001000110011: color_data = 12'b110011001100;
		14'b01001000110100: color_data = 12'b110011001100;
		14'b01001000110101: color_data = 12'b110011001100;
		14'b01001000110110: color_data = 12'b110011001100;
		14'b01001000110111: color_data = 12'b110011001100;
		14'b01001000111000: color_data = 12'b110011001100;
		14'b01001000111001: color_data = 12'b110011001100;
		14'b01001000111010: color_data = 12'b110011001100;
		14'b01001000111011: color_data = 12'b110011001100;
		14'b01001000111100: color_data = 12'b110011001100;
		14'b01001000111101: color_data = 12'b110011001100;
		14'b01001000111110: color_data = 12'b110011001100;
		14'b01001000111111: color_data = 12'b110011001100;
		14'b01001001000000: color_data = 12'b110011001100;
		14'b01001001000001: color_data = 12'b110011001100;
		14'b01001001000010: color_data = 12'b110011001100;
		14'b01001001000011: color_data = 12'b110011001100;
		14'b01001001000100: color_data = 12'b110011001100;
		14'b01001001000101: color_data = 12'b110011001100;
		14'b01001001000110: color_data = 12'b110011001100;
		14'b01001001000111: color_data = 12'b110011001100;
		14'b01001001001000: color_data = 12'b110011001100;
		14'b01001001001001: color_data = 12'b110011001100;
		14'b01001001001010: color_data = 12'b110011001100;
		14'b01001001001011: color_data = 12'b011101110111;
		14'b01001010010111: color_data = 12'b000000000000;
		14'b01001010011000: color_data = 12'b111000010010;
		14'b01001010011001: color_data = 12'b111000010010;
		14'b01001010011010: color_data = 12'b111000010010;
		14'b01001010011011: color_data = 12'b111000010010;
		14'b01001010011100: color_data = 12'b111000010010;
		14'b01001010011101: color_data = 12'b111000010010;
		14'b01001010011110: color_data = 12'b111000010010;
		14'b01001010011111: color_data = 12'b111000010010;
		14'b01001010100000: color_data = 12'b111000010010;
		14'b01001010100001: color_data = 12'b111000010010;
		14'b01001010100010: color_data = 12'b111000010010;
		14'b01001010100011: color_data = 12'b111000010010;
		14'b01001010100100: color_data = 12'b111000010010;
		14'b01001010100101: color_data = 12'b111000010010;
		14'b01001010100110: color_data = 12'b111000010010;
		14'b01001010100111: color_data = 12'b111000010010;
		14'b01001010101000: color_data = 12'b111000010010;
		14'b01001010101001: color_data = 12'b011101110111;
		14'b01001010101010: color_data = 12'b110011001100;
		14'b01001010101011: color_data = 12'b110011001100;
		14'b01001010101100: color_data = 12'b110011001100;
		14'b01001010101101: color_data = 12'b110011001100;
		14'b01001010101110: color_data = 12'b110011001100;
		14'b01001010101111: color_data = 12'b110011001100;
		14'b01001010110000: color_data = 12'b110011001100;
		14'b01001010110001: color_data = 12'b110011001100;
		14'b01001010110010: color_data = 12'b110011001100;
		14'b01001010110011: color_data = 12'b110011001100;
		14'b01001010110100: color_data = 12'b110011001100;
		14'b01001010110101: color_data = 12'b110011001100;
		14'b01001010110110: color_data = 12'b110011001100;
		14'b01001010110111: color_data = 12'b110011001100;
		14'b01001010111000: color_data = 12'b110011001100;
		14'b01001010111001: color_data = 12'b110011001100;
		14'b01001010111010: color_data = 12'b110011001100;
		14'b01001010111011: color_data = 12'b110011001100;
		14'b01001010111100: color_data = 12'b110011001100;
		14'b01001010111101: color_data = 12'b110011001100;
		14'b01001010111110: color_data = 12'b110011001100;
		14'b01001010111111: color_data = 12'b110011001100;
		14'b01001011000000: color_data = 12'b110011001100;
		14'b01001011000001: color_data = 12'b110011001100;
		14'b01001011000010: color_data = 12'b110011001100;
		14'b01001011000011: color_data = 12'b110011001100;
		14'b01001011000100: color_data = 12'b110011001100;
		14'b01001011000101: color_data = 12'b110011001100;
		14'b01001011000110: color_data = 12'b110011001100;
		14'b01001011000111: color_data = 12'b110011001100;
		14'b01001011001000: color_data = 12'b110011001100;
		14'b01001011001001: color_data = 12'b110011001100;
		14'b01001011001010: color_data = 12'b110011001100;
		14'b01001011001011: color_data = 12'b011101110111;
		14'b01001100010111: color_data = 12'b000000000000;
		14'b01001100011000: color_data = 12'b111000010010;
		14'b01001100011001: color_data = 12'b111000010010;
		14'b01001100011010: color_data = 12'b111000010010;
		14'b01001100011011: color_data = 12'b111000010010;
		14'b01001100011100: color_data = 12'b111000010010;
		14'b01001100011101: color_data = 12'b111000010010;
		14'b01001100011110: color_data = 12'b111000010010;
		14'b01001100011111: color_data = 12'b111000010010;
		14'b01001100100000: color_data = 12'b111000010010;
		14'b01001100100001: color_data = 12'b111000010010;
		14'b01001100100010: color_data = 12'b111000010010;
		14'b01001100100011: color_data = 12'b111000010010;
		14'b01001100100100: color_data = 12'b111000010010;
		14'b01001100100101: color_data = 12'b111000010010;
		14'b01001100100110: color_data = 12'b111000010010;
		14'b01001100100111: color_data = 12'b111000010010;
		14'b01001100101000: color_data = 12'b111000010010;
		14'b01001100101001: color_data = 12'b011101110111;
		14'b01001100101010: color_data = 12'b110011001100;
		14'b01001100101011: color_data = 12'b110011001100;
		14'b01001100101100: color_data = 12'b110011001100;
		14'b01001100101101: color_data = 12'b110011001100;
		14'b01001100101110: color_data = 12'b110011001100;
		14'b01001100101111: color_data = 12'b110011001100;
		14'b01001100110000: color_data = 12'b110011001100;
		14'b01001100110001: color_data = 12'b110011001100;
		14'b01001100110010: color_data = 12'b110011001100;
		14'b01001100110011: color_data = 12'b110011001100;
		14'b01001100110100: color_data = 12'b110011001100;
		14'b01001100110101: color_data = 12'b110011001100;
		14'b01001100110110: color_data = 12'b110011001100;
		14'b01001100110111: color_data = 12'b110011001100;
		14'b01001100111000: color_data = 12'b110011001100;
		14'b01001100111001: color_data = 12'b110011001100;
		14'b01001100111010: color_data = 12'b110011001100;
		14'b01001100111011: color_data = 12'b110011001100;
		14'b01001100111100: color_data = 12'b110011001100;
		14'b01001100111101: color_data = 12'b110011001100;
		14'b01001100111110: color_data = 12'b110011001100;
		14'b01001100111111: color_data = 12'b110011001100;
		14'b01001101000000: color_data = 12'b110011001100;
		14'b01001101000001: color_data = 12'b110011001100;
		14'b01001101000010: color_data = 12'b110011001100;
		14'b01001101000011: color_data = 12'b110011001100;
		14'b01001101000100: color_data = 12'b110011001100;
		14'b01001101000101: color_data = 12'b110011001100;
		14'b01001101000110: color_data = 12'b110011001100;
		14'b01001101000111: color_data = 12'b110011001100;
		14'b01001101001000: color_data = 12'b110011001100;
		14'b01001101001001: color_data = 12'b110011001100;
		14'b01001101001010: color_data = 12'b110011001100;
		14'b01001101001011: color_data = 12'b011101110111;
		14'b01001110010111: color_data = 12'b000000000000;
		14'b01001110011000: color_data = 12'b111000010010;
		14'b01001110011001: color_data = 12'b111000010010;
		14'b01001110011010: color_data = 12'b111000010010;
		14'b01001110011011: color_data = 12'b111000010010;
		14'b01001110011100: color_data = 12'b111000010010;
		14'b01001110011101: color_data = 12'b111000010010;
		14'b01001110011110: color_data = 12'b111000010010;
		14'b01001110011111: color_data = 12'b111000010010;
		14'b01001110100000: color_data = 12'b111000010010;
		14'b01001110100001: color_data = 12'b111000010010;
		14'b01001110100010: color_data = 12'b111000010010;
		14'b01001110100011: color_data = 12'b111000010010;
		14'b01001110100100: color_data = 12'b111000010010;
		14'b01001110100101: color_data = 12'b111000010010;
		14'b01001110100110: color_data = 12'b111000010010;
		14'b01001110100111: color_data = 12'b111000010010;
		14'b01001110101000: color_data = 12'b111000010010;
		14'b01001110101001: color_data = 12'b011101110111;
		14'b01001110101010: color_data = 12'b110011001100;
		14'b01001110101011: color_data = 12'b110011001100;
		14'b01001110101100: color_data = 12'b110011001100;
		14'b01001110101101: color_data = 12'b110011001100;
		14'b01001110101110: color_data = 12'b110011001100;
		14'b01001110101111: color_data = 12'b110011001100;
		14'b01001110110000: color_data = 12'b110011001100;
		14'b01001110110001: color_data = 12'b110011001100;
		14'b01001110110010: color_data = 12'b110011001100;
		14'b01001110110011: color_data = 12'b110011001100;
		14'b01001110110100: color_data = 12'b110011001100;
		14'b01001110110101: color_data = 12'b110011001100;
		14'b01001110110110: color_data = 12'b110011001100;
		14'b01001110110111: color_data = 12'b110011001100;
		14'b01001110111000: color_data = 12'b110011001100;
		14'b01001110111001: color_data = 12'b110011001100;
		14'b01001110111010: color_data = 12'b110011001100;
		14'b01001110111011: color_data = 12'b110011001100;
		14'b01001110111100: color_data = 12'b110011001100;
		14'b01001110111101: color_data = 12'b110011001100;
		14'b01001110111110: color_data = 12'b110011001100;
		14'b01001110111111: color_data = 12'b110011001100;
		14'b01001111000000: color_data = 12'b110011001100;
		14'b01001111000001: color_data = 12'b110011001100;
		14'b01001111000010: color_data = 12'b110011001100;
		14'b01001111000011: color_data = 12'b110011001100;
		14'b01001111000100: color_data = 12'b110011001100;
		14'b01001111000101: color_data = 12'b110011001100;
		14'b01001111000110: color_data = 12'b110011001100;
		14'b01001111000111: color_data = 12'b110011001100;
		14'b01001111001000: color_data = 12'b110011001100;
		14'b01001111001001: color_data = 12'b110011001100;
		14'b01001111001010: color_data = 12'b110011001100;
		14'b01001111001011: color_data = 12'b011101110111;
		14'b01010000010111: color_data = 12'b000000000000;
		14'b01010000011000: color_data = 12'b111000010010;
		14'b01010000011001: color_data = 12'b111000010010;
		14'b01010000011010: color_data = 12'b111000010010;
		14'b01010000011011: color_data = 12'b111000010010;
		14'b01010000011100: color_data = 12'b111000010010;
		14'b01010000011101: color_data = 12'b111000010010;
		14'b01010000011110: color_data = 12'b111000010010;
		14'b01010000011111: color_data = 12'b111000010010;
		14'b01010000100000: color_data = 12'b111000010010;
		14'b01010000100001: color_data = 12'b111000010010;
		14'b01010000100010: color_data = 12'b111000010010;
		14'b01010000100011: color_data = 12'b111000010010;
		14'b01010000100100: color_data = 12'b111000010010;
		14'b01010000100101: color_data = 12'b111000010010;
		14'b01010000100110: color_data = 12'b111000010010;
		14'b01010000100111: color_data = 12'b111000010010;
		14'b01010000101000: color_data = 12'b111000010010;
		14'b01010000101001: color_data = 12'b011101110111;
		14'b01010000101010: color_data = 12'b110011001100;
		14'b01010000101011: color_data = 12'b110011001100;
		14'b01010000101100: color_data = 12'b110011001100;
		14'b01010000101101: color_data = 12'b110011001100;
		14'b01010000101110: color_data = 12'b110011001100;
		14'b01010000101111: color_data = 12'b110011001100;
		14'b01010000110000: color_data = 12'b110011001100;
		14'b01010000110001: color_data = 12'b110011001100;
		14'b01010000110010: color_data = 12'b110011001100;
		14'b01010000110011: color_data = 12'b110011001100;
		14'b01010000110100: color_data = 12'b110011001100;
		14'b01010000110101: color_data = 12'b110011001100;
		14'b01010000110110: color_data = 12'b110011001100;
		14'b01010000110111: color_data = 12'b110011001100;
		14'b01010000111000: color_data = 12'b110011001100;
		14'b01010000111001: color_data = 12'b110011001100;
		14'b01010000111010: color_data = 12'b110011001100;
		14'b01010000111011: color_data = 12'b110011001100;
		14'b01010000111100: color_data = 12'b110011001100;
		14'b01010000111101: color_data = 12'b110011001100;
		14'b01010000111110: color_data = 12'b110011001100;
		14'b01010000111111: color_data = 12'b110011001100;
		14'b01010001000000: color_data = 12'b110011001100;
		14'b01010001000001: color_data = 12'b110011001100;
		14'b01010001000010: color_data = 12'b110011001100;
		14'b01010001000011: color_data = 12'b110011001100;
		14'b01010001000100: color_data = 12'b110011001100;
		14'b01010001000101: color_data = 12'b110011001100;
		14'b01010001000110: color_data = 12'b110011001100;
		14'b01010001000111: color_data = 12'b110011001100;
		14'b01010001001000: color_data = 12'b110011001100;
		14'b01010001001001: color_data = 12'b110011001100;
		14'b01010001001010: color_data = 12'b110011001100;
		14'b01010001001011: color_data = 12'b011101110111;
		14'b01010010010111: color_data = 12'b000000000000;
		14'b01010010011000: color_data = 12'b111000010010;
		14'b01010010011001: color_data = 12'b111000010010;
		14'b01010010011010: color_data = 12'b111000010010;
		14'b01010010011011: color_data = 12'b111000010010;
		14'b01010010011100: color_data = 12'b111000010010;
		14'b01010010011101: color_data = 12'b111000010010;
		14'b01010010011110: color_data = 12'b111000010010;
		14'b01010010011111: color_data = 12'b111000010010;
		14'b01010010100000: color_data = 12'b111000010010;
		14'b01010010100001: color_data = 12'b111000010010;
		14'b01010010100010: color_data = 12'b111000010010;
		14'b01010010100011: color_data = 12'b111000010010;
		14'b01010010100100: color_data = 12'b111000010010;
		14'b01010010100101: color_data = 12'b111000010010;
		14'b01010010100110: color_data = 12'b111000010010;
		14'b01010010100111: color_data = 12'b111000010010;
		14'b01010010101000: color_data = 12'b111000010010;
		14'b01010010101001: color_data = 12'b011101110111;
		14'b01010010101010: color_data = 12'b110011001100;
		14'b01010010101011: color_data = 12'b110011001100;
		14'b01010010101100: color_data = 12'b110011001100;
		14'b01010010101101: color_data = 12'b110011001100;
		14'b01010010101110: color_data = 12'b110011001100;
		14'b01010010101111: color_data = 12'b110011001100;
		14'b01010010110000: color_data = 12'b110011001100;
		14'b01010010110001: color_data = 12'b110011001100;
		14'b01010010110010: color_data = 12'b110011001100;
		14'b01010010110011: color_data = 12'b110011001100;
		14'b01010010110100: color_data = 12'b110011001100;
		14'b01010010110101: color_data = 12'b110011001100;
		14'b01010010110110: color_data = 12'b110011001100;
		14'b01010010110111: color_data = 12'b110011001100;
		14'b01010010111000: color_data = 12'b110011001100;
		14'b01010010111001: color_data = 12'b110011001100;
		14'b01010010111010: color_data = 12'b110011001100;
		14'b01010010111011: color_data = 12'b110011001100;
		14'b01010010111100: color_data = 12'b110011001100;
		14'b01010010111101: color_data = 12'b110011001100;
		14'b01010010111110: color_data = 12'b110011001100;
		14'b01010010111111: color_data = 12'b110011001100;
		14'b01010011000000: color_data = 12'b110011001100;
		14'b01010011000001: color_data = 12'b110011001100;
		14'b01010011000010: color_data = 12'b110011001100;
		14'b01010011000011: color_data = 12'b110011001100;
		14'b01010011000100: color_data = 12'b110011001100;
		14'b01010011000101: color_data = 12'b110011001100;
		14'b01010011000110: color_data = 12'b110011001100;
		14'b01010011000111: color_data = 12'b110011001100;
		14'b01010011001000: color_data = 12'b110011001100;
		14'b01010011001001: color_data = 12'b110011001100;
		14'b01010011001010: color_data = 12'b110011001100;
		14'b01010011001011: color_data = 12'b011101110111;
		14'b01010100010111: color_data = 12'b000000000000;
		14'b01010100011000: color_data = 12'b111000010010;
		14'b01010100011001: color_data = 12'b111000010010;
		14'b01010100011010: color_data = 12'b111000010010;
		14'b01010100011011: color_data = 12'b111000010010;
		14'b01010100011100: color_data = 12'b111000010010;
		14'b01010100011101: color_data = 12'b111000010010;
		14'b01010100011110: color_data = 12'b111000010010;
		14'b01010100011111: color_data = 12'b111000010010;
		14'b01010100100000: color_data = 12'b111000010010;
		14'b01010100100001: color_data = 12'b111000010010;
		14'b01010100100010: color_data = 12'b111000010010;
		14'b01010100100011: color_data = 12'b111000010010;
		14'b01010100100100: color_data = 12'b111000010010;
		14'b01010100100101: color_data = 12'b111000010010;
		14'b01010100100110: color_data = 12'b111000010010;
		14'b01010100100111: color_data = 12'b111000010010;
		14'b01010100101000: color_data = 12'b111000010010;
		14'b01010100101001: color_data = 12'b011101110111;
		14'b01010100101010: color_data = 12'b110011001100;
		14'b01010100101011: color_data = 12'b110011001100;
		14'b01010100101100: color_data = 12'b110011001100;
		14'b01010100101101: color_data = 12'b110011001100;
		14'b01010100101110: color_data = 12'b110011001100;
		14'b01010100101111: color_data = 12'b110011001100;
		14'b01010100110000: color_data = 12'b110011001100;
		14'b01010100110001: color_data = 12'b110011001100;
		14'b01010100110010: color_data = 12'b110011001100;
		14'b01010100110011: color_data = 12'b110011001100;
		14'b01010100110100: color_data = 12'b110011001100;
		14'b01010100110101: color_data = 12'b110011001100;
		14'b01010100110110: color_data = 12'b110011001100;
		14'b01010100110111: color_data = 12'b110011001100;
		14'b01010100111000: color_data = 12'b110011001100;
		14'b01010100111001: color_data = 12'b110011001100;
		14'b01010100111010: color_data = 12'b110011001100;
		14'b01010100111011: color_data = 12'b110011001100;
		14'b01010100111100: color_data = 12'b110011001100;
		14'b01010100111101: color_data = 12'b110011001100;
		14'b01010100111110: color_data = 12'b110011001100;
		14'b01010100111111: color_data = 12'b110011001100;
		14'b01010101000000: color_data = 12'b110011001100;
		14'b01010101000001: color_data = 12'b110011001100;
		14'b01010101000010: color_data = 12'b110011001100;
		14'b01010101000011: color_data = 12'b110011001100;
		14'b01010101000100: color_data = 12'b110011001100;
		14'b01010101000101: color_data = 12'b110011001100;
		14'b01010101000110: color_data = 12'b110011001100;
		14'b01010101000111: color_data = 12'b110011001100;
		14'b01010101001000: color_data = 12'b110011001100;
		14'b01010101001001: color_data = 12'b110011001100;
		14'b01010101001010: color_data = 12'b110011001100;
		14'b01010101001011: color_data = 12'b011101110111;
		14'b01010110010111: color_data = 12'b000000000000;
		14'b01010110011000: color_data = 12'b111000010010;
		14'b01010110011001: color_data = 12'b111000010010;
		14'b01010110011010: color_data = 12'b111000010010;
		14'b01010110011011: color_data = 12'b111000010010;
		14'b01010110011100: color_data = 12'b111000010010;
		14'b01010110011101: color_data = 12'b111000010010;
		14'b01010110011110: color_data = 12'b111000010010;
		14'b01010110011111: color_data = 12'b111000010010;
		14'b01010110100000: color_data = 12'b111000010010;
		14'b01010110100001: color_data = 12'b111000010010;
		14'b01010110100010: color_data = 12'b111000010010;
		14'b01010110100011: color_data = 12'b111000010010;
		14'b01010110100100: color_data = 12'b111000010010;
		14'b01010110100101: color_data = 12'b111000010010;
		14'b01010110100110: color_data = 12'b111000010010;
		14'b01010110100111: color_data = 12'b111000010010;
		14'b01010110101000: color_data = 12'b111000010010;
		14'b01010110101001: color_data = 12'b011101110111;
		14'b01010110101010: color_data = 12'b110011001100;
		14'b01010110101011: color_data = 12'b110011001100;
		14'b01010110101100: color_data = 12'b110011001100;
		14'b01010110101101: color_data = 12'b110011001100;
		14'b01010110101110: color_data = 12'b110011001100;
		14'b01010110101111: color_data = 12'b110011001100;
		14'b01010110110000: color_data = 12'b110011001100;
		14'b01010110110001: color_data = 12'b110011001100;
		14'b01010110110010: color_data = 12'b110011001100;
		14'b01010110110011: color_data = 12'b110011001100;
		14'b01010110110100: color_data = 12'b110011001100;
		14'b01010110110101: color_data = 12'b110011001100;
		14'b01010110110110: color_data = 12'b110011001100;
		14'b01010110110111: color_data = 12'b110011001100;
		14'b01010110111000: color_data = 12'b110011001100;
		14'b01010110111001: color_data = 12'b110011001100;
		14'b01010110111010: color_data = 12'b110011001100;
		14'b01010110111011: color_data = 12'b110011001100;
		14'b01010110111100: color_data = 12'b110011001100;
		14'b01010110111101: color_data = 12'b110011001100;
		14'b01010110111110: color_data = 12'b110011001100;
		14'b01010110111111: color_data = 12'b110011001100;
		14'b01010111000000: color_data = 12'b110011001100;
		14'b01010111000001: color_data = 12'b110011001100;
		14'b01010111000010: color_data = 12'b110011001100;
		14'b01010111000011: color_data = 12'b110011001100;
		14'b01010111000100: color_data = 12'b110011001100;
		14'b01010111000101: color_data = 12'b110011001100;
		14'b01010111000110: color_data = 12'b110011001100;
		14'b01010111000111: color_data = 12'b110011001100;
		14'b01010111001000: color_data = 12'b110011001100;
		14'b01010111001001: color_data = 12'b110011001100;
		14'b01010111001010: color_data = 12'b110011001100;
		14'b01010111001011: color_data = 12'b011101110111;
		14'b01011000010111: color_data = 12'b000000000000;
		14'b01011000011000: color_data = 12'b111000010010;
		14'b01011000011001: color_data = 12'b111000010010;
		14'b01011000011010: color_data = 12'b111000010010;
		14'b01011000011011: color_data = 12'b111000010010;
		14'b01011000011100: color_data = 12'b111000010010;
		14'b01011000011101: color_data = 12'b111000010010;
		14'b01011000011110: color_data = 12'b111000010010;
		14'b01011000011111: color_data = 12'b111000010010;
		14'b01011000100000: color_data = 12'b111000010010;
		14'b01011000100001: color_data = 12'b111000010010;
		14'b01011000100010: color_data = 12'b111000010010;
		14'b01011000100011: color_data = 12'b111000010010;
		14'b01011000100100: color_data = 12'b111000010010;
		14'b01011000100101: color_data = 12'b111000010010;
		14'b01011000100110: color_data = 12'b111000010010;
		14'b01011000100111: color_data = 12'b111000010010;
		14'b01011000101000: color_data = 12'b111000010010;
		14'b01011000101001: color_data = 12'b011101110111;
		14'b01011000101010: color_data = 12'b110011001100;
		14'b01011000101011: color_data = 12'b110011001100;
		14'b01011000101100: color_data = 12'b110011001100;
		14'b01011000101101: color_data = 12'b110011001100;
		14'b01011000101110: color_data = 12'b110011001100;
		14'b01011000101111: color_data = 12'b110011001100;
		14'b01011000110000: color_data = 12'b110011001100;
		14'b01011000110001: color_data = 12'b110011001100;
		14'b01011000110010: color_data = 12'b110011001100;
		14'b01011000110011: color_data = 12'b110011001100;
		14'b01011000110100: color_data = 12'b110011001100;
		14'b01011000110101: color_data = 12'b110011001100;
		14'b01011000110110: color_data = 12'b110011001100;
		14'b01011000110111: color_data = 12'b110011001100;
		14'b01011000111000: color_data = 12'b110011001100;
		14'b01011000111001: color_data = 12'b110011001100;
		14'b01011000111010: color_data = 12'b110011001100;
		14'b01011000111011: color_data = 12'b110011001100;
		14'b01011000111100: color_data = 12'b110011001100;
		14'b01011000111101: color_data = 12'b110011001100;
		14'b01011000111110: color_data = 12'b110011001100;
		14'b01011000111111: color_data = 12'b110011001100;
		14'b01011001000000: color_data = 12'b110011001100;
		14'b01011001000001: color_data = 12'b110011001100;
		14'b01011001000010: color_data = 12'b110011001100;
		14'b01011001000011: color_data = 12'b110011001100;
		14'b01011001000100: color_data = 12'b110011001100;
		14'b01011001000101: color_data = 12'b110011001100;
		14'b01011001000110: color_data = 12'b110011001100;
		14'b01011001000111: color_data = 12'b110011001100;
		14'b01011001001000: color_data = 12'b110011001100;
		14'b01011001001001: color_data = 12'b110011001100;
		14'b01011001001010: color_data = 12'b110011001100;
		14'b01011001001011: color_data = 12'b011101110111;
		14'b01011010010111: color_data = 12'b000000000000;
		14'b01011010011000: color_data = 12'b111000010010;
		14'b01011010011001: color_data = 12'b111000010010;
		14'b01011010011010: color_data = 12'b111000010010;
		14'b01011010011011: color_data = 12'b111000010010;
		14'b01011010011100: color_data = 12'b111000010010;
		14'b01011010011101: color_data = 12'b111000010010;
		14'b01011010011110: color_data = 12'b111000010010;
		14'b01011010011111: color_data = 12'b111000010010;
		14'b01011010100000: color_data = 12'b111000010010;
		14'b01011010100001: color_data = 12'b111000010010;
		14'b01011010100010: color_data = 12'b111000010010;
		14'b01011010100011: color_data = 12'b111000010010;
		14'b01011010100100: color_data = 12'b111000010010;
		14'b01011010100101: color_data = 12'b111000010010;
		14'b01011010100110: color_data = 12'b111000010010;
		14'b01011010100111: color_data = 12'b111000010010;
		14'b01011010101000: color_data = 12'b111000010010;
		14'b01011010101001: color_data = 12'b011101110111;
		14'b01011010101010: color_data = 12'b110011001100;
		14'b01011010101011: color_data = 12'b110011001100;
		14'b01011010101100: color_data = 12'b011101110111;
		14'b01011010101101: color_data = 12'b110011001100;
		14'b01011010101110: color_data = 12'b110011001100;
		14'b01011010101111: color_data = 12'b110011001100;
		14'b01011010110000: color_data = 12'b110011001100;
		14'b01011010110001: color_data = 12'b110011001100;
		14'b01011010110010: color_data = 12'b110011001100;
		14'b01011010110011: color_data = 12'b110011001100;
		14'b01011010110100: color_data = 12'b110011001100;
		14'b01011010110101: color_data = 12'b110011001100;
		14'b01011010110110: color_data = 12'b110011001100;
		14'b01011010110111: color_data = 12'b110011001100;
		14'b01011010111000: color_data = 12'b110011001100;
		14'b01011010111001: color_data = 12'b110011001100;
		14'b01011010111010: color_data = 12'b110011001100;
		14'b01011010111011: color_data = 12'b110011001100;
		14'b01011010111100: color_data = 12'b110011001100;
		14'b01011010111101: color_data = 12'b110011001100;
		14'b01011010111110: color_data = 12'b110011001100;
		14'b01011010111111: color_data = 12'b110011001100;
		14'b01011011000000: color_data = 12'b110011001100;
		14'b01011011000001: color_data = 12'b110011001100;
		14'b01011011000010: color_data = 12'b110011001100;
		14'b01011011000011: color_data = 12'b110011001100;
		14'b01011011000100: color_data = 12'b110011001100;
		14'b01011011000101: color_data = 12'b110011001100;
		14'b01011011000110: color_data = 12'b110011001100;
		14'b01011011000111: color_data = 12'b110011001100;
		14'b01011011001000: color_data = 12'b110011001100;
		14'b01011011001001: color_data = 12'b011101110111;
		14'b01011011001010: color_data = 12'b110011001100;
		14'b01011011001011: color_data = 12'b011101110111;
		14'b01011100010111: color_data = 12'b000000000000;
		14'b01011100011000: color_data = 12'b111000010010;
		14'b01011100011001: color_data = 12'b111000010010;
		14'b01011100011010: color_data = 12'b111000010010;
		14'b01011100011011: color_data = 12'b111000010010;
		14'b01011100011100: color_data = 12'b111000010010;
		14'b01011100011101: color_data = 12'b111000010010;
		14'b01011100011110: color_data = 12'b111000010010;
		14'b01011100011111: color_data = 12'b111000010010;
		14'b01011100100000: color_data = 12'b111000010010;
		14'b01011100100001: color_data = 12'b111000010010;
		14'b01011100100010: color_data = 12'b111000010010;
		14'b01011100100011: color_data = 12'b111000010010;
		14'b01011100100100: color_data = 12'b111000010010;
		14'b01011100100101: color_data = 12'b111000010010;
		14'b01011100100110: color_data = 12'b111000010010;
		14'b01011100100111: color_data = 12'b111000010010;
		14'b01011100101000: color_data = 12'b111000010010;
		14'b01011100101001: color_data = 12'b011101110111;
		14'b01011100101010: color_data = 12'b110011001100;
		14'b01011100101011: color_data = 12'b110011001100;
		14'b01011100101100: color_data = 12'b110011001100;
		14'b01011100101101: color_data = 12'b110011001100;
		14'b01011100101110: color_data = 12'b110011001100;
		14'b01011100101111: color_data = 12'b110011001100;
		14'b01011100110000: color_data = 12'b110011001100;
		14'b01011100110001: color_data = 12'b110011001100;
		14'b01011100110010: color_data = 12'b110011001100;
		14'b01011100110011: color_data = 12'b110011001100;
		14'b01011100110100: color_data = 12'b110011001100;
		14'b01011100110101: color_data = 12'b110011001100;
		14'b01011100110110: color_data = 12'b110011001100;
		14'b01011100110111: color_data = 12'b110011001100;
		14'b01011100111000: color_data = 12'b110011001100;
		14'b01011100111001: color_data = 12'b110011001100;
		14'b01011100111010: color_data = 12'b110011001100;
		14'b01011100111011: color_data = 12'b110011001100;
		14'b01011100111100: color_data = 12'b110011001100;
		14'b01011100111101: color_data = 12'b110011001100;
		14'b01011100111110: color_data = 12'b110011001100;
		14'b01011100111111: color_data = 12'b110011001100;
		14'b01011101000000: color_data = 12'b110011001100;
		14'b01011101000001: color_data = 12'b110011001100;
		14'b01011101000010: color_data = 12'b110011001100;
		14'b01011101000011: color_data = 12'b110011001100;
		14'b01011101000100: color_data = 12'b110011001100;
		14'b01011101000101: color_data = 12'b110011001100;
		14'b01011101000110: color_data = 12'b110011001100;
		14'b01011101000111: color_data = 12'b110011001100;
		14'b01011101001000: color_data = 12'b110011001100;
		14'b01011101001001: color_data = 12'b110011001100;
		14'b01011101001010: color_data = 12'b110011001100;
		14'b01011101001011: color_data = 12'b011101110111;
		14'b01011110010111: color_data = 12'b000000000000;
		14'b01011110011000: color_data = 12'b111000010010;
		14'b01011110011001: color_data = 12'b111000010010;
		14'b01011110011010: color_data = 12'b111000010010;
		14'b01011110011011: color_data = 12'b111000010010;
		14'b01011110011100: color_data = 12'b111000010010;
		14'b01011110011101: color_data = 12'b111000010010;
		14'b01011110011110: color_data = 12'b111000010010;
		14'b01011110011111: color_data = 12'b111000010010;
		14'b01011110100000: color_data = 12'b111000010010;
		14'b01011110100001: color_data = 12'b111000010010;
		14'b01011110100010: color_data = 12'b111000010010;
		14'b01011110100011: color_data = 12'b111000010010;
		14'b01011110100100: color_data = 12'b111000010010;
		14'b01011110100101: color_data = 12'b111000010010;
		14'b01011110100110: color_data = 12'b111000010010;
		14'b01011110100111: color_data = 12'b111000010010;
		14'b01011110101000: color_data = 12'b111000010010;
		14'b01011110101001: color_data = 12'b111000010010;
		14'b01011110101010: color_data = 12'b011101110111;
		14'b01011110101011: color_data = 12'b011101110111;
		14'b01011110101100: color_data = 12'b110011001100;
		14'b01011110101101: color_data = 12'b110011001100;
		14'b01011110101110: color_data = 12'b110011001100;
		14'b01011110101111: color_data = 12'b110011001100;
		14'b01011110110000: color_data = 12'b110011001100;
		14'b01011110110001: color_data = 12'b110011001100;
		14'b01011110110010: color_data = 12'b110011001100;
		14'b01011110110011: color_data = 12'b110011001100;
		14'b01011110110100: color_data = 12'b110011001100;
		14'b01011110110101: color_data = 12'b110011001100;
		14'b01011110110110: color_data = 12'b110011001100;
		14'b01011110110111: color_data = 12'b110011001100;
		14'b01011110111000: color_data = 12'b110011001100;
		14'b01011110111001: color_data = 12'b110011001100;
		14'b01011110111010: color_data = 12'b110011001100;
		14'b01011110111011: color_data = 12'b110011001100;
		14'b01011110111100: color_data = 12'b110011001100;
		14'b01011110111101: color_data = 12'b110011001100;
		14'b01011110111110: color_data = 12'b110011001100;
		14'b01011110111111: color_data = 12'b110011001100;
		14'b01011111000000: color_data = 12'b110011001100;
		14'b01011111000001: color_data = 12'b110011001100;
		14'b01011111000010: color_data = 12'b110011001100;
		14'b01011111000011: color_data = 12'b110011001100;
		14'b01011111000100: color_data = 12'b110011001100;
		14'b01011111000101: color_data = 12'b110011001100;
		14'b01011111000110: color_data = 12'b110011001100;
		14'b01011111000111: color_data = 12'b110011001100;
		14'b01011111001000: color_data = 12'b110011001100;
		14'b01011111001001: color_data = 12'b011101110111;
		14'b01011111001010: color_data = 12'b011101110111;
		14'b01100000010111: color_data = 12'b000000000000;
		14'b01100000011000: color_data = 12'b111000010010;
		14'b01100000011001: color_data = 12'b111000010010;
		14'b01100000011010: color_data = 12'b111000010010;
		14'b01100000011011: color_data = 12'b111000010010;
		14'b01100000011100: color_data = 12'b111000010010;
		14'b01100000011101: color_data = 12'b111000010010;
		14'b01100000011110: color_data = 12'b111000010010;
		14'b01100000011111: color_data = 12'b111000010010;
		14'b01100000100000: color_data = 12'b111000010010;
		14'b01100000100001: color_data = 12'b111000010010;
		14'b01100000100010: color_data = 12'b111000010010;
		14'b01100000100011: color_data = 12'b111000010010;
		14'b01100000100100: color_data = 12'b111000010010;
		14'b01100000100101: color_data = 12'b111000010010;
		14'b01100000100110: color_data = 12'b111000010010;
		14'b01100000100111: color_data = 12'b111000010010;
		14'b01100000101000: color_data = 12'b111000010010;
		14'b01100000101001: color_data = 12'b111000010010;
		14'b01100000101010: color_data = 12'b111000010010;
		14'b01100000101011: color_data = 12'b111000010010;
		14'b01100000101100: color_data = 12'b011101110111;
		14'b01100000101101: color_data = 12'b011101110111;
		14'b01100000101110: color_data = 12'b110011001100;
		14'b01100000101111: color_data = 12'b110011001100;
		14'b01100000110000: color_data = 12'b110011001100;
		14'b01100000110001: color_data = 12'b110011001100;
		14'b01100000110010: color_data = 12'b110011001100;
		14'b01100000110011: color_data = 12'b110011001100;
		14'b01100000110100: color_data = 12'b110011001100;
		14'b01100000110101: color_data = 12'b110011001100;
		14'b01100000110110: color_data = 12'b110011001100;
		14'b01100000110111: color_data = 12'b110011001100;
		14'b01100000111000: color_data = 12'b110011001100;
		14'b01100000111001: color_data = 12'b110011001100;
		14'b01100000111010: color_data = 12'b110011001100;
		14'b01100000111011: color_data = 12'b110011001100;
		14'b01100000111100: color_data = 12'b110011001100;
		14'b01100000111101: color_data = 12'b110011001100;
		14'b01100000111110: color_data = 12'b110011001100;
		14'b01100000111111: color_data = 12'b110011001100;
		14'b01100001000000: color_data = 12'b110011001100;
		14'b01100001000001: color_data = 12'b110011001100;
		14'b01100001000010: color_data = 12'b110011001100;
		14'b01100001000011: color_data = 12'b110011001100;
		14'b01100001000100: color_data = 12'b110011001100;
		14'b01100001000101: color_data = 12'b110011001100;
		14'b01100001000110: color_data = 12'b110011001100;
		14'b01100001000111: color_data = 12'b011101110111;
		14'b01100001001000: color_data = 12'b011101110111;
		14'b01100010010111: color_data = 12'b000000000000;
		14'b01100010011000: color_data = 12'b111000010010;
		14'b01100010011001: color_data = 12'b111000010010;
		14'b01100010011010: color_data = 12'b111000010010;
		14'b01100010011011: color_data = 12'b111000010010;
		14'b01100010011100: color_data = 12'b111000010010;
		14'b01100010011101: color_data = 12'b111000010010;
		14'b01100010011110: color_data = 12'b111000010010;
		14'b01100010011111: color_data = 12'b111000010010;
		14'b01100010100000: color_data = 12'b111000010010;
		14'b01100010100001: color_data = 12'b111000010010;
		14'b01100010100010: color_data = 12'b111000010010;
		14'b01100010100011: color_data = 12'b111000010010;
		14'b01100010100100: color_data = 12'b111000010010;
		14'b01100010100101: color_data = 12'b111000010010;
		14'b01100010100110: color_data = 12'b111000010010;
		14'b01100010100111: color_data = 12'b111000010010;
		14'b01100010101000: color_data = 12'b111000010010;
		14'b01100010101001: color_data = 12'b111000010010;
		14'b01100010101010: color_data = 12'b111000010010;
		14'b01100010101011: color_data = 12'b111000010010;
		14'b01100010101100: color_data = 12'b111000010010;
		14'b01100010101101: color_data = 12'b111000010010;
		14'b01100010101110: color_data = 12'b011101110111;
		14'b01100010101111: color_data = 12'b110011001100;
		14'b01100010110000: color_data = 12'b110011001100;
		14'b01100010110001: color_data = 12'b110011001100;
		14'b01100010110010: color_data = 12'b110011001100;
		14'b01100010110011: color_data = 12'b110011001100;
		14'b01100010110100: color_data = 12'b110011001100;
		14'b01100010110101: color_data = 12'b110011001100;
		14'b01100010110110: color_data = 12'b110011001100;
		14'b01100010110111: color_data = 12'b110011001100;
		14'b01100010111000: color_data = 12'b110011001100;
		14'b01100010111001: color_data = 12'b110011001100;
		14'b01100010111010: color_data = 12'b110011001100;
		14'b01100010111011: color_data = 12'b110011001100;
		14'b01100010111100: color_data = 12'b110011001100;
		14'b01100010111101: color_data = 12'b110011001100;
		14'b01100010111110: color_data = 12'b110011001100;
		14'b01100010111111: color_data = 12'b110011001100;
		14'b01100011000000: color_data = 12'b110011001100;
		14'b01100011000001: color_data = 12'b110011001100;
		14'b01100011000010: color_data = 12'b110011001100;
		14'b01100011000011: color_data = 12'b110011001100;
		14'b01100011000100: color_data = 12'b110011001100;
		14'b01100011000101: color_data = 12'b110011001100;
		14'b01100011000110: color_data = 12'b011101110111;
		14'b01100100010111: color_data = 12'b000000000000;
		14'b01100100011000: color_data = 12'b111000010010;
		14'b01100100011001: color_data = 12'b111000010010;
		14'b01100100011010: color_data = 12'b111000010010;
		14'b01100100011011: color_data = 12'b111000010010;
		14'b01100100011100: color_data = 12'b111000010010;
		14'b01100100011101: color_data = 12'b111000010010;
		14'b01100100011110: color_data = 12'b111000010010;
		14'b01100100011111: color_data = 12'b111000010010;
		14'b01100100100000: color_data = 12'b111000010010;
		14'b01100100100001: color_data = 12'b111000010010;
		14'b01100100100010: color_data = 12'b111000010010;
		14'b01100100100011: color_data = 12'b111000010010;
		14'b01100100100100: color_data = 12'b111000010010;
		14'b01100100100101: color_data = 12'b111000010010;
		14'b01100100100110: color_data = 12'b111000010010;
		14'b01100100100111: color_data = 12'b111000010010;
		14'b01100100101000: color_data = 12'b111000010010;
		14'b01100100101001: color_data = 12'b111000010010;
		14'b01100100101010: color_data = 12'b111000010010;
		14'b01100100101011: color_data = 12'b111000010010;
		14'b01100100101100: color_data = 12'b111000010010;
		14'b01100100101101: color_data = 12'b111000010010;
		14'b01100100101110: color_data = 12'b111000010010;
		14'b01100100101111: color_data = 12'b011101110111;
		14'b01100100110000: color_data = 12'b011101110111;
		14'b01100100110001: color_data = 12'b110011001100;
		14'b01100100110010: color_data = 12'b110011001100;
		14'b01100100110011: color_data = 12'b110011001100;
		14'b01100100110100: color_data = 12'b110011001100;
		14'b01100100110101: color_data = 12'b110011001100;
		14'b01100100110110: color_data = 12'b110011001100;
		14'b01100100110111: color_data = 12'b110011001100;
		14'b01100100111000: color_data = 12'b110011001100;
		14'b01100100111001: color_data = 12'b110011001100;
		14'b01100100111010: color_data = 12'b110011001100;
		14'b01100100111011: color_data = 12'b110011001100;
		14'b01100100111100: color_data = 12'b110011001100;
		14'b01100100111101: color_data = 12'b110011001100;
		14'b01100100111110: color_data = 12'b110011001100;
		14'b01100100111111: color_data = 12'b110011001100;
		14'b01100101000000: color_data = 12'b110011001100;
		14'b01100101000001: color_data = 12'b110011001100;
		14'b01100101000010: color_data = 12'b110011001100;
		14'b01100101000011: color_data = 12'b110011001100;
		14'b01100101000100: color_data = 12'b011101110111;
		14'b01100101000101: color_data = 12'b011101110111;
		14'b01100110010111: color_data = 12'b000000000000;
		14'b01100110011000: color_data = 12'b111000010010;
		14'b01100110011001: color_data = 12'b111000010010;
		14'b01100110011010: color_data = 12'b111000010010;
		14'b01100110011011: color_data = 12'b111000010010;
		14'b01100110011100: color_data = 12'b111000010010;
		14'b01100110011101: color_data = 12'b111000010010;
		14'b01100110011110: color_data = 12'b111000010010;
		14'b01100110011111: color_data = 12'b111000010010;
		14'b01100110100000: color_data = 12'b111000010010;
		14'b01100110100001: color_data = 12'b111000010010;
		14'b01100110100010: color_data = 12'b111000010010;
		14'b01100110100011: color_data = 12'b111000010010;
		14'b01100110100100: color_data = 12'b111000010010;
		14'b01100110100101: color_data = 12'b111000010010;
		14'b01100110100110: color_data = 12'b111000010010;
		14'b01100110100111: color_data = 12'b111000010010;
		14'b01100110101000: color_data = 12'b111000010010;
		14'b01100110101001: color_data = 12'b111000010010;
		14'b01100110101010: color_data = 12'b111000010010;
		14'b01100110101011: color_data = 12'b111000010010;
		14'b01100110101100: color_data = 12'b111000010010;
		14'b01100110101101: color_data = 12'b111000010010;
		14'b01100110101110: color_data = 12'b111000010010;
		14'b01100110101111: color_data = 12'b111000010010;
		14'b01100110110000: color_data = 12'b000000000000;
		14'b01100110110001: color_data = 12'b011101110111;
		14'b01100110110010: color_data = 12'b011101110111;
		14'b01100110110011: color_data = 12'b110011001100;
		14'b01100110110100: color_data = 12'b110011001100;
		14'b01100110110101: color_data = 12'b110011001100;
		14'b01100110110110: color_data = 12'b110011001100;
		14'b01100110110111: color_data = 12'b110011001100;
		14'b01100110111000: color_data = 12'b110011001100;
		14'b01100110111001: color_data = 12'b110011001100;
		14'b01100110111010: color_data = 12'b110011001100;
		14'b01100110111011: color_data = 12'b110011001100;
		14'b01100110111100: color_data = 12'b110011001100;
		14'b01100110111101: color_data = 12'b110011001100;
		14'b01100110111110: color_data = 12'b110011001100;
		14'b01100110111111: color_data = 12'b110011001100;
		14'b01100111000000: color_data = 12'b110011001100;
		14'b01100111000001: color_data = 12'b110011001100;
		14'b01100111000010: color_data = 12'b011101110111;
		14'b01100111000011: color_data = 12'b011101110111;
		14'b01101000010111: color_data = 12'b000000000000;
		14'b01101000011000: color_data = 12'b111000010010;
		14'b01101000011001: color_data = 12'b111000010010;
		14'b01101000011010: color_data = 12'b111000010010;
		14'b01101000011011: color_data = 12'b111000010010;
		14'b01101000011100: color_data = 12'b111000010010;
		14'b01101000011101: color_data = 12'b111000010010;
		14'b01101000011110: color_data = 12'b111000010010;
		14'b01101000011111: color_data = 12'b111000010010;
		14'b01101000100000: color_data = 12'b111000010010;
		14'b01101000100001: color_data = 12'b111000010010;
		14'b01101000100010: color_data = 12'b111000010010;
		14'b01101000100011: color_data = 12'b111000010010;
		14'b01101000100100: color_data = 12'b111000010010;
		14'b01101000100101: color_data = 12'b111000010010;
		14'b01101000100110: color_data = 12'b111000010010;
		14'b01101000100111: color_data = 12'b111000010010;
		14'b01101000101000: color_data = 12'b111000010010;
		14'b01101000101001: color_data = 12'b111000010010;
		14'b01101000101010: color_data = 12'b111000010010;
		14'b01101000101011: color_data = 12'b111000010010;
		14'b01101000101100: color_data = 12'b111000010010;
		14'b01101000101101: color_data = 12'b111000010010;
		14'b01101000101110: color_data = 12'b111000010010;
		14'b01101000101111: color_data = 12'b111000010010;
		14'b01101000110000: color_data = 12'b000000000000;
		14'b01101000110011: color_data = 12'b011101110111;
		14'b01101000110100: color_data = 12'b011101110111;
		14'b01101000110101: color_data = 12'b110011001100;
		14'b01101000110110: color_data = 12'b110011001100;
		14'b01101000110111: color_data = 12'b110011001100;
		14'b01101000111000: color_data = 12'b110011001100;
		14'b01101000111001: color_data = 12'b110011001100;
		14'b01101000111010: color_data = 12'b110011001100;
		14'b01101000111011: color_data = 12'b110011001100;
		14'b01101000111100: color_data = 12'b110011001100;
		14'b01101000111101: color_data = 12'b110011001100;
		14'b01101000111110: color_data = 12'b110011001100;
		14'b01101000111111: color_data = 12'b110011001100;
		14'b01101001000000: color_data = 12'b011101110111;
		14'b01101001000001: color_data = 12'b011101110111;
		14'b01101010010111: color_data = 12'b000000000000;
		14'b01101010011000: color_data = 12'b111000010010;
		14'b01101010011001: color_data = 12'b111000010010;
		14'b01101010011010: color_data = 12'b111000010010;
		14'b01101010011011: color_data = 12'b111000010010;
		14'b01101010011100: color_data = 12'b111000010010;
		14'b01101010011101: color_data = 12'b111000010010;
		14'b01101010011110: color_data = 12'b111000010010;
		14'b01101010011111: color_data = 12'b111000010010;
		14'b01101010100000: color_data = 12'b111000010010;
		14'b01101010100001: color_data = 12'b111000010010;
		14'b01101010100010: color_data = 12'b111000010010;
		14'b01101010100011: color_data = 12'b111000010010;
		14'b01101010100100: color_data = 12'b111000010010;
		14'b01101010100101: color_data = 12'b111000010010;
		14'b01101010100110: color_data = 12'b111000010010;
		14'b01101010100111: color_data = 12'b111000010010;
		14'b01101010101000: color_data = 12'b111000010010;
		14'b01101010101001: color_data = 12'b111000010010;
		14'b01101010101010: color_data = 12'b111000010010;
		14'b01101010101011: color_data = 12'b111000010010;
		14'b01101010101100: color_data = 12'b111000010010;
		14'b01101010101101: color_data = 12'b111000010010;
		14'b01101010101110: color_data = 12'b111000010010;
		14'b01101010101111: color_data = 12'b111000010010;
		14'b01101010110000: color_data = 12'b000000000000;
		14'b01101010110101: color_data = 12'b011101110111;
		14'b01101010110110: color_data = 12'b110011001100;
		14'b01101010110111: color_data = 12'b110011001100;
		14'b01101010111000: color_data = 12'b110011001100;
		14'b01101010111001: color_data = 12'b110011001100;
		14'b01101010111010: color_data = 12'b011101110111;
		14'b01101010111011: color_data = 12'b110011001100;
		14'b01101010111100: color_data = 12'b110011001100;
		14'b01101010111101: color_data = 12'b110011001100;
		14'b01101010111110: color_data = 12'b110011001100;
		14'b01101010111111: color_data = 12'b011101110111;
		14'b01101100010111: color_data = 12'b000000000000;
		14'b01101100011000: color_data = 12'b111000010010;
		14'b01101100011001: color_data = 12'b111000010010;
		14'b01101100011010: color_data = 12'b111000010010;
		14'b01101100011011: color_data = 12'b111000010010;
		14'b01101100011100: color_data = 12'b111000010010;
		14'b01101100011101: color_data = 12'b111000010010;
		14'b01101100011110: color_data = 12'b111000010010;
		14'b01101100011111: color_data = 12'b111000010010;
		14'b01101100100000: color_data = 12'b111000010010;
		14'b01101100100001: color_data = 12'b111000010010;
		14'b01101100100010: color_data = 12'b111000010010;
		14'b01101100100011: color_data = 12'b111000010010;
		14'b01101100100100: color_data = 12'b111000010010;
		14'b01101100100101: color_data = 12'b111000010010;
		14'b01101100100110: color_data = 12'b111000010010;
		14'b01101100100111: color_data = 12'b111000010010;
		14'b01101100101000: color_data = 12'b111000010010;
		14'b01101100101001: color_data = 12'b111000010010;
		14'b01101100101010: color_data = 12'b111000010010;
		14'b01101100101011: color_data = 12'b111000010010;
		14'b01101100101100: color_data = 12'b111000010010;
		14'b01101100101101: color_data = 12'b111000010010;
		14'b01101100101110: color_data = 12'b111000010010;
		14'b01101100101111: color_data = 12'b111000010010;
		14'b01101100110000: color_data = 12'b000000000000;
		14'b01101100110110: color_data = 12'b011101110111;
		14'b01101100110111: color_data = 12'b011101110111;
		14'b01101100111000: color_data = 12'b110011001100;
		14'b01101100111001: color_data = 12'b110011001100;
		14'b01101100111010: color_data = 12'b110011001100;
		14'b01101100111011: color_data = 12'b110011001100;
		14'b01101100111100: color_data = 12'b110011001100;
		14'b01101100111101: color_data = 12'b011101110111;
		14'b01101100111110: color_data = 12'b011101110111;
		14'b01101110010111: color_data = 12'b000000000000;
		14'b01101110011000: color_data = 12'b111000010010;
		14'b01101110011001: color_data = 12'b111000010010;
		14'b01101110011010: color_data = 12'b111000010010;
		14'b01101110011011: color_data = 12'b111000010010;
		14'b01101110011100: color_data = 12'b111000010010;
		14'b01101110011101: color_data = 12'b111000010010;
		14'b01101110011110: color_data = 12'b111000010010;
		14'b01101110011111: color_data = 12'b111000010010;
		14'b01101110100000: color_data = 12'b111000010010;
		14'b01101110100001: color_data = 12'b111000010010;
		14'b01101110100010: color_data = 12'b111000010010;
		14'b01101110100011: color_data = 12'b111000010010;
		14'b01101110100100: color_data = 12'b111000010010;
		14'b01101110100101: color_data = 12'b111000010010;
		14'b01101110100110: color_data = 12'b111000010010;
		14'b01101110100111: color_data = 12'b111000010010;
		14'b01101110101000: color_data = 12'b111000010010;
		14'b01101110101001: color_data = 12'b111000010010;
		14'b01101110101010: color_data = 12'b111000010010;
		14'b01101110101011: color_data = 12'b111000010010;
		14'b01101110101100: color_data = 12'b111000010010;
		14'b01101110101101: color_data = 12'b111000010010;
		14'b01101110101110: color_data = 12'b111000010010;
		14'b01101110101111: color_data = 12'b111000010010;
		14'b01101110110000: color_data = 12'b000000000000;
		14'b01101110111000: color_data = 12'b011101110111;
		14'b01101110111001: color_data = 12'b011101110111;
		14'b01101110111010: color_data = 12'b110011001100;
		14'b01101110111011: color_data = 12'b011101110111;
		14'b01101110111100: color_data = 12'b011101110111;
		14'b01110000010111: color_data = 12'b000000000000;
		14'b01110000011000: color_data = 12'b111000010010;
		14'b01110000011001: color_data = 12'b111000010010;
		14'b01110000011010: color_data = 12'b111000010010;
		14'b01110000011011: color_data = 12'b111000010010;
		14'b01110000011100: color_data = 12'b111000010010;
		14'b01110000011101: color_data = 12'b111000010010;
		14'b01110000011110: color_data = 12'b111000010010;
		14'b01110000011111: color_data = 12'b111000010010;
		14'b01110000100000: color_data = 12'b111000010010;
		14'b01110000100001: color_data = 12'b111000010010;
		14'b01110000100010: color_data = 12'b111000010010;
		14'b01110000100011: color_data = 12'b111000010010;
		14'b01110000100100: color_data = 12'b111000010010;
		14'b01110000100101: color_data = 12'b111000010010;
		14'b01110000100110: color_data = 12'b111000010010;
		14'b01110000100111: color_data = 12'b111000010010;
		14'b01110000101000: color_data = 12'b111000010010;
		14'b01110000101001: color_data = 12'b111000010010;
		14'b01110000101010: color_data = 12'b111000010010;
		14'b01110000101011: color_data = 12'b111000010010;
		14'b01110000101100: color_data = 12'b111000010010;
		14'b01110000101101: color_data = 12'b111000010010;
		14'b01110000101110: color_data = 12'b111000010010;
		14'b01110000101111: color_data = 12'b111000010010;
		14'b01110000110000: color_data = 12'b000000000000;
		14'b01110000111010: color_data = 12'b011101110111;
		14'b01110010010111: color_data = 12'b000000000000;
		14'b01110010011000: color_data = 12'b111000010010;
		14'b01110010011001: color_data = 12'b111000010010;
		14'b01110010011010: color_data = 12'b111000010010;
		14'b01110010011011: color_data = 12'b111000010010;
		14'b01110010011100: color_data = 12'b111000010010;
		14'b01110010011101: color_data = 12'b111000010010;
		14'b01110010011110: color_data = 12'b111000010010;
		14'b01110010011111: color_data = 12'b111000010010;
		14'b01110010100000: color_data = 12'b111000010010;
		14'b01110010100001: color_data = 12'b111000010010;
		14'b01110010100010: color_data = 12'b111000010010;
		14'b01110010100011: color_data = 12'b111000010010;
		14'b01110010100100: color_data = 12'b111000010010;
		14'b01110010100101: color_data = 12'b111000010010;
		14'b01110010100110: color_data = 12'b111000010010;
		14'b01110010100111: color_data = 12'b111000010010;
		14'b01110010101000: color_data = 12'b111000010010;
		14'b01110010101001: color_data = 12'b111000010010;
		14'b01110010101010: color_data = 12'b111000010010;
		14'b01110010101011: color_data = 12'b111000010010;
		14'b01110010101100: color_data = 12'b111000010010;
		14'b01110010101101: color_data = 12'b111000010010;
		14'b01110010101110: color_data = 12'b111000010010;
		14'b01110010101111: color_data = 12'b111000010010;
		14'b01110010110000: color_data = 12'b000000000000;
		14'b01110100010111: color_data = 12'b000000000000;
		14'b01110100011000: color_data = 12'b111000010010;
		14'b01110100011001: color_data = 12'b111000010010;
		14'b01110100011010: color_data = 12'b111000010010;
		14'b01110100011011: color_data = 12'b111000010010;
		14'b01110100011100: color_data = 12'b111000010010;
		14'b01110100011101: color_data = 12'b111000010010;
		14'b01110100011110: color_data = 12'b111000010010;
		14'b01110100011111: color_data = 12'b111000010010;
		14'b01110100100000: color_data = 12'b111000010010;
		14'b01110100100001: color_data = 12'b111000010010;
		14'b01110100100010: color_data = 12'b111000010010;
		14'b01110100100011: color_data = 12'b111000010010;
		14'b01110100100100: color_data = 12'b111000010010;
		14'b01110100100101: color_data = 12'b111000010010;
		14'b01110100100110: color_data = 12'b111000010010;
		14'b01110100100111: color_data = 12'b111000010010;
		14'b01110100101000: color_data = 12'b111000010010;
		14'b01110100101001: color_data = 12'b111000010010;
		14'b01110100101010: color_data = 12'b111000010010;
		14'b01110100101011: color_data = 12'b111000010010;
		14'b01110100101100: color_data = 12'b111000010010;
		14'b01110100101101: color_data = 12'b111000010010;
		14'b01110100101110: color_data = 12'b111000010010;
		14'b01110100101111: color_data = 12'b111000010010;
		14'b01110100110000: color_data = 12'b000000000000;
		14'b01110110010111: color_data = 12'b000000000000;
		14'b01110110011000: color_data = 12'b111000010010;
		14'b01110110011001: color_data = 12'b111000010010;
		14'b01110110011010: color_data = 12'b111000010010;
		14'b01110110011011: color_data = 12'b111000010010;
		14'b01110110011100: color_data = 12'b111000010010;
		14'b01110110011101: color_data = 12'b111000010010;
		14'b01110110011110: color_data = 12'b111000010010;
		14'b01110110011111: color_data = 12'b111000010010;
		14'b01110110100000: color_data = 12'b111000010010;
		14'b01110110100001: color_data = 12'b111000010010;
		14'b01110110100010: color_data = 12'b111000010010;
		14'b01110110100011: color_data = 12'b111000010010;
		14'b01110110100100: color_data = 12'b111000010010;
		14'b01110110100101: color_data = 12'b111000010010;
		14'b01110110100110: color_data = 12'b111000010010;
		14'b01110110100111: color_data = 12'b111000010010;
		14'b01110110101000: color_data = 12'b111000010010;
		14'b01110110101001: color_data = 12'b111000010010;
		14'b01110110101010: color_data = 12'b111000010010;
		14'b01110110101011: color_data = 12'b111000010010;
		14'b01110110101100: color_data = 12'b111000010010;
		14'b01110110101101: color_data = 12'b111000010010;
		14'b01110110101110: color_data = 12'b111000010010;
		14'b01110110101111: color_data = 12'b111000010010;
		14'b01110110110000: color_data = 12'b000000000000;
		14'b01111000010111: color_data = 12'b000000000000;
		14'b01111000011000: color_data = 12'b111000010010;
		14'b01111000011001: color_data = 12'b111000010010;
		14'b01111000011010: color_data = 12'b111000010010;
		14'b01111000011011: color_data = 12'b111000010010;
		14'b01111000011100: color_data = 12'b111000010010;
		14'b01111000011101: color_data = 12'b111000010010;
		14'b01111000011110: color_data = 12'b111000010010;
		14'b01111000011111: color_data = 12'b111000010010;
		14'b01111000100000: color_data = 12'b111000010010;
		14'b01111000100001: color_data = 12'b111000010010;
		14'b01111000100010: color_data = 12'b111000010010;
		14'b01111000100011: color_data = 12'b111000010010;
		14'b01111000100100: color_data = 12'b111000010010;
		14'b01111000100101: color_data = 12'b111000010010;
		14'b01111000100110: color_data = 12'b111000010010;
		14'b01111000100111: color_data = 12'b111000010010;
		14'b01111000101000: color_data = 12'b111000010010;
		14'b01111000101001: color_data = 12'b111000010010;
		14'b01111000101010: color_data = 12'b111000010010;
		14'b01111000101011: color_data = 12'b111000010010;
		14'b01111000101100: color_data = 12'b111000010010;
		14'b01111000101101: color_data = 12'b111000010010;
		14'b01111000101110: color_data = 12'b111000010010;
		14'b01111000101111: color_data = 12'b111000010010;
		14'b01111000110000: color_data = 12'b000000000000;
		14'b01111010010111: color_data = 12'b000000000000;
		14'b01111010011000: color_data = 12'b001101001100;
		14'b01111010011001: color_data = 12'b001101001100;
		14'b01111010011010: color_data = 12'b001101001100;
		14'b01111010011011: color_data = 12'b001101001100;
		14'b01111010011100: color_data = 12'b001101001100;
		14'b01111010011101: color_data = 12'b001101001100;
		14'b01111010011110: color_data = 12'b001101001100;
		14'b01111010011111: color_data = 12'b001101001100;
		14'b01111010100000: color_data = 12'b001101001100;
		14'b01111010100001: color_data = 12'b001101001100;
		14'b01111010100010: color_data = 12'b001101001100;
		14'b01111010100011: color_data = 12'b001101001100;
		14'b01111010100100: color_data = 12'b001101001100;
		14'b01111010100101: color_data = 12'b001101001100;
		14'b01111010100110: color_data = 12'b001101001100;
		14'b01111010100111: color_data = 12'b001101001100;
		14'b01111010101000: color_data = 12'b001101001100;
		14'b01111010101001: color_data = 12'b001101001100;
		14'b01111010101010: color_data = 12'b001101001100;
		14'b01111010101011: color_data = 12'b001101001100;
		14'b01111010101100: color_data = 12'b001101001100;
		14'b01111010101101: color_data = 12'b001101001100;
		14'b01111010101110: color_data = 12'b001101001100;
		14'b01111010101111: color_data = 12'b001101001100;
		14'b01111010110000: color_data = 12'b000000000000;
		14'b01111100010111: color_data = 12'b000000000000;
		14'b01111100011000: color_data = 12'b001101001100;
		14'b01111100011001: color_data = 12'b001101001100;
		14'b01111100011010: color_data = 12'b001101001100;
		14'b01111100011011: color_data = 12'b001101001100;
		14'b01111100011100: color_data = 12'b001101001100;
		14'b01111100011101: color_data = 12'b001101001100;
		14'b01111100011110: color_data = 12'b001101001100;
		14'b01111100011111: color_data = 12'b001101001100;
		14'b01111100100000: color_data = 12'b001101001100;
		14'b01111100100001: color_data = 12'b001101001100;
		14'b01111100100010: color_data = 12'b001101001100;
		14'b01111100100011: color_data = 12'b001101001100;
		14'b01111100100100: color_data = 12'b001101001100;
		14'b01111100100101: color_data = 12'b001101001100;
		14'b01111100100110: color_data = 12'b001101001100;
		14'b01111100100111: color_data = 12'b001101001100;
		14'b01111100101000: color_data = 12'b001101001100;
		14'b01111100101001: color_data = 12'b001101001100;
		14'b01111100101010: color_data = 12'b001101001100;
		14'b01111100101011: color_data = 12'b001101001100;
		14'b01111100101100: color_data = 12'b001101001100;
		14'b01111100101101: color_data = 12'b001101001100;
		14'b01111100101110: color_data = 12'b001101001100;
		14'b01111100101111: color_data = 12'b001101001100;
		14'b01111100110000: color_data = 12'b000000000000;
		14'b01111110010111: color_data = 12'b000000000000;
		14'b01111110011000: color_data = 12'b001101001100;
		14'b01111110011001: color_data = 12'b001101001100;
		14'b01111110011010: color_data = 12'b001101001100;
		14'b01111110011011: color_data = 12'b001101001100;
		14'b01111110011100: color_data = 12'b001101001100;
		14'b01111110011101: color_data = 12'b001101001100;
		14'b01111110011110: color_data = 12'b001101001100;
		14'b01111110011111: color_data = 12'b001101001100;
		14'b01111110100000: color_data = 12'b001101001100;
		14'b01111110100001: color_data = 12'b001101001100;
		14'b01111110100010: color_data = 12'b001101001100;
		14'b01111110100011: color_data = 12'b001101001100;
		14'b01111110100100: color_data = 12'b001101001100;
		14'b01111110100101: color_data = 12'b001101001100;
		14'b01111110100110: color_data = 12'b001101001100;
		14'b01111110100111: color_data = 12'b001101001100;
		14'b01111110101000: color_data = 12'b001101001100;
		14'b01111110101001: color_data = 12'b001101001100;
		14'b01111110101010: color_data = 12'b001101001100;
		14'b01111110101011: color_data = 12'b001101001100;
		14'b01111110101100: color_data = 12'b001101001100;
		14'b01111110101101: color_data = 12'b001101001100;
		14'b01111110101110: color_data = 12'b001101001100;
		14'b01111110101111: color_data = 12'b001101001100;
		14'b01111110110000: color_data = 12'b000000000000;
		14'b10000000010111: color_data = 12'b000000000000;
		14'b10000000011000: color_data = 12'b001101001100;
		14'b10000000011001: color_data = 12'b001101001100;
		14'b10000000011010: color_data = 12'b001101001100;
		14'b10000000011011: color_data = 12'b001101001100;
		14'b10000000011100: color_data = 12'b001101001100;
		14'b10000000011101: color_data = 12'b001101001100;
		14'b10000000011110: color_data = 12'b001101001100;
		14'b10000000011111: color_data = 12'b001101001100;
		14'b10000000100000: color_data = 12'b001101001100;
		14'b10000000100001: color_data = 12'b001101001100;
		14'b10000000100010: color_data = 12'b001101001100;
		14'b10000000100011: color_data = 12'b001101001100;
		14'b10000000100100: color_data = 12'b001101001100;
		14'b10000000100101: color_data = 12'b001101001100;
		14'b10000000100110: color_data = 12'b001101001100;
		14'b10000000100111: color_data = 12'b001101001100;
		14'b10000000101000: color_data = 12'b001101001100;
		14'b10000000101001: color_data = 12'b001101001100;
		14'b10000000101010: color_data = 12'b001101001100;
		14'b10000000101011: color_data = 12'b001101001100;
		14'b10000000101100: color_data = 12'b001101001100;
		14'b10000000101101: color_data = 12'b001101001100;
		14'b10000000101110: color_data = 12'b001101001100;
		14'b10000000101111: color_data = 12'b001101001100;
		14'b10000000110000: color_data = 12'b000000000000;
		14'b10000010010111: color_data = 12'b000000000000;
		14'b10000010011000: color_data = 12'b001101001100;
		14'b10000010011001: color_data = 12'b001101001100;
		14'b10000010011010: color_data = 12'b001101001100;
		14'b10000010011011: color_data = 12'b001101001100;
		14'b10000010011100: color_data = 12'b001101001100;
		14'b10000010011101: color_data = 12'b001101001100;
		14'b10000010011110: color_data = 12'b001101001100;
		14'b10000010011111: color_data = 12'b001101001100;
		14'b10000010100000: color_data = 12'b001101001100;
		14'b10000010100001: color_data = 12'b001101001100;
		14'b10000010100010: color_data = 12'b001101001100;
		14'b10000010100011: color_data = 12'b001101001100;
		14'b10000010100100: color_data = 12'b001101001100;
		14'b10000010100101: color_data = 12'b001101001100;
		14'b10000010100110: color_data = 12'b001101001100;
		14'b10000010100111: color_data = 12'b001101001100;
		14'b10000010101000: color_data = 12'b001101001100;
		14'b10000010101001: color_data = 12'b001101001100;
		14'b10000010101010: color_data = 12'b001101001100;
		14'b10000010101011: color_data = 12'b001101001100;
		14'b10000010101100: color_data = 12'b001101001100;
		14'b10000010101101: color_data = 12'b001101001100;
		14'b10000010101110: color_data = 12'b001101001100;
		14'b10000010101111: color_data = 12'b001101001100;
		14'b10000010110000: color_data = 12'b000000000000;
		14'b10000100010111: color_data = 12'b000000000000;
		14'b10000100011000: color_data = 12'b001101001100;
		14'b10000100011001: color_data = 12'b001101001100;
		14'b10000100011010: color_data = 12'b001101001100;
		14'b10000100011011: color_data = 12'b001101001100;
		14'b10000100011100: color_data = 12'b001101001100;
		14'b10000100011101: color_data = 12'b001101001100;
		14'b10000100011110: color_data = 12'b000000000000;
		14'b10000100011111: color_data = 12'b000000000000;
		14'b10000100100000: color_data = 12'b000000000000;
		14'b10000100100001: color_data = 12'b000000000000;
		14'b10000100100010: color_data = 12'b000000000000;
		14'b10000100100011: color_data = 12'b000000000000;
		14'b10000100100100: color_data = 12'b000000000000;
		14'b10000100100101: color_data = 12'b000000000000;
		14'b10000100100110: color_data = 12'b000000000000;
		14'b10000100100111: color_data = 12'b000000000000;
		14'b10000100101000: color_data = 12'b000000000000;
		14'b10000100101001: color_data = 12'b000000000000;
		14'b10000100101010: color_data = 12'b001101001100;
		14'b10000100101011: color_data = 12'b001101001100;
		14'b10000100101100: color_data = 12'b001101001100;
		14'b10000100101101: color_data = 12'b001101001100;
		14'b10000100101110: color_data = 12'b001101001100;
		14'b10000100101111: color_data = 12'b001101001100;
		14'b10000100110000: color_data = 12'b000000000000;
		14'b10000110010111: color_data = 12'b000000000000;
		14'b10000110011000: color_data = 12'b001101001100;
		14'b10000110011001: color_data = 12'b001101001100;
		14'b10000110011010: color_data = 12'b001101001100;
		14'b10000110011011: color_data = 12'b001101001100;
		14'b10000110011100: color_data = 12'b001101001100;
		14'b10000110011101: color_data = 12'b001101001100;
		14'b10000110011110: color_data = 12'b000000000000;
		14'b10000110101001: color_data = 12'b000000000000;
		14'b10000110101010: color_data = 12'b001101001100;
		14'b10000110101011: color_data = 12'b001101001100;
		14'b10000110101100: color_data = 12'b001101001100;
		14'b10000110101101: color_data = 12'b001101001100;
		14'b10000110101110: color_data = 12'b001101001100;
		14'b10000110101111: color_data = 12'b001101001100;
		14'b10000110110000: color_data = 12'b000000000000;
		14'b10001000010111: color_data = 12'b000000000000;
		14'b10001000011000: color_data = 12'b001101001100;
		14'b10001000011001: color_data = 12'b001101001100;
		14'b10001000011010: color_data = 12'b001101001100;
		14'b10001000011011: color_data = 12'b001101001100;
		14'b10001000011100: color_data = 12'b001101001100;
		14'b10001000011101: color_data = 12'b001101001100;
		14'b10001000011110: color_data = 12'b000000000000;
		14'b10001000101001: color_data = 12'b000000000000;
		14'b10001000101010: color_data = 12'b001101001100;
		14'b10001000101011: color_data = 12'b001101001100;
		14'b10001000101100: color_data = 12'b001101001100;
		14'b10001000101101: color_data = 12'b001101001100;
		14'b10001000101110: color_data = 12'b001101001100;
		14'b10001000101111: color_data = 12'b001101001100;
		14'b10001000110000: color_data = 12'b000000000000;
		14'b10001010010111: color_data = 12'b000000000000;
		14'b10001010011000: color_data = 12'b001101001100;
		14'b10001010011001: color_data = 12'b001101001100;
		14'b10001010011010: color_data = 12'b001101001100;
		14'b10001010011011: color_data = 12'b001101001100;
		14'b10001010011100: color_data = 12'b001101001100;
		14'b10001010011101: color_data = 12'b001101001100;
		14'b10001010011110: color_data = 12'b000000000000;
		14'b10001010101001: color_data = 12'b000000000000;
		14'b10001010101010: color_data = 12'b001101001100;
		14'b10001010101011: color_data = 12'b001101001100;
		14'b10001010101100: color_data = 12'b001101001100;
		14'b10001010101101: color_data = 12'b001101001100;
		14'b10001010101110: color_data = 12'b001101001100;
		14'b10001010101111: color_data = 12'b001101001100;
		14'b10001010110000: color_data = 12'b000000000000;
		14'b10001100010111: color_data = 12'b000000000000;
		14'b10001100011000: color_data = 12'b001101001100;
		14'b10001100011001: color_data = 12'b001101001100;
		14'b10001100011010: color_data = 12'b001101001100;
		14'b10001100011011: color_data = 12'b001101001100;
		14'b10001100011100: color_data = 12'b001101001100;
		14'b10001100011101: color_data = 12'b001101001100;
		14'b10001100011110: color_data = 12'b000000000000;
		14'b10001100101001: color_data = 12'b000000000000;
		14'b10001100101010: color_data = 12'b001101001100;
		14'b10001100101011: color_data = 12'b001101001100;
		14'b10001100101100: color_data = 12'b001101001100;
		14'b10001100101101: color_data = 12'b001101001100;
		14'b10001100101110: color_data = 12'b001101001100;
		14'b10001100101111: color_data = 12'b001101001100;
		14'b10001100110000: color_data = 12'b000000000000;
		14'b10001110010111: color_data = 12'b000000000000;
		14'b10001110011000: color_data = 12'b001101001100;
		14'b10001110011001: color_data = 12'b001101001100;
		14'b10001110011010: color_data = 12'b001101001100;
		14'b10001110011011: color_data = 12'b001101001100;
		14'b10001110011100: color_data = 12'b001101001100;
		14'b10001110011101: color_data = 12'b001101001100;
		14'b10001110011110: color_data = 12'b000000000000;
		14'b10001110101001: color_data = 12'b000000000000;
		14'b10001110101010: color_data = 12'b001101001100;
		14'b10001110101011: color_data = 12'b001101001100;
		14'b10001110101100: color_data = 12'b001101001100;
		14'b10001110101101: color_data = 12'b001101001100;
		14'b10001110101110: color_data = 12'b001101001100;
		14'b10001110101111: color_data = 12'b001101001100;
		14'b10001110110000: color_data = 12'b000000000000;
		14'b10010000010111: color_data = 12'b000000000000;
		14'b10010000011000: color_data = 12'b001101001100;
		14'b10010000011001: color_data = 12'b001101001100;
		14'b10010000011010: color_data = 12'b001101001100;
		14'b10010000011011: color_data = 12'b001101001100;
		14'b10010000011100: color_data = 12'b001101001100;
		14'b10010000011101: color_data = 12'b001101001100;
		14'b10010000011110: color_data = 12'b000000000000;
		14'b10010000101001: color_data = 12'b000000000000;
		14'b10010000101010: color_data = 12'b001101001100;
		14'b10010000101011: color_data = 12'b001101001100;
		14'b10010000101100: color_data = 12'b001101001100;
		14'b10010000101101: color_data = 12'b001101001100;
		14'b10010000101110: color_data = 12'b001101001100;
		14'b10010000101111: color_data = 12'b001101001100;
		14'b10010000110000: color_data = 12'b000000000000;
		14'b10010010010111: color_data = 12'b000000000000;
		14'b10010010011000: color_data = 12'b001101001100;
		14'b10010010011001: color_data = 12'b001101001100;
		14'b10010010011010: color_data = 12'b001101001100;
		14'b10010010011011: color_data = 12'b001101001100;
		14'b10010010011100: color_data = 12'b001101001100;
		14'b10010010011101: color_data = 12'b001101001100;
		14'b10010010011110: color_data = 12'b000000000000;
		14'b10010010101001: color_data = 12'b000000000000;
		14'b10010010101010: color_data = 12'b001101001100;
		14'b10010010101011: color_data = 12'b001101001100;
		14'b10010010101100: color_data = 12'b001101001100;
		14'b10010010101101: color_data = 12'b001101001100;
		14'b10010010101110: color_data = 12'b001101001100;
		14'b10010010101111: color_data = 12'b001101001100;
		14'b10010010110000: color_data = 12'b000000000000;
		14'b10010100010111: color_data = 12'b000000000000;
		14'b10010100011000: color_data = 12'b001101001100;
		14'b10010100011001: color_data = 12'b001101001100;
		14'b10010100011010: color_data = 12'b001101001100;
		14'b10010100011011: color_data = 12'b001101001100;
		14'b10010100011100: color_data = 12'b001101001100;
		14'b10010100011101: color_data = 12'b001101001100;
		14'b10010100011110: color_data = 12'b000000000000;
		14'b10010100101001: color_data = 12'b000000000000;
		14'b10010100101010: color_data = 12'b001101001100;
		14'b10010100101011: color_data = 12'b001101001100;
		14'b10010100101100: color_data = 12'b001101001100;
		14'b10010100101101: color_data = 12'b001101001100;
		14'b10010100101110: color_data = 12'b001101001100;
		14'b10010100101111: color_data = 12'b001101001100;
		14'b10010100110000: color_data = 12'b000000000000;
		14'b10010110010111: color_data = 12'b000000000000;
		14'b10010110011000: color_data = 12'b001101001100;
		14'b10010110011001: color_data = 12'b001101001100;
		14'b10010110011010: color_data = 12'b001101001100;
		14'b10010110011011: color_data = 12'b001101001100;
		14'b10010110011100: color_data = 12'b001101001100;
		14'b10010110011101: color_data = 12'b001101001100;
		14'b10010110011110: color_data = 12'b000000000000;
		14'b10010110101001: color_data = 12'b000000000000;
		14'b10010110101010: color_data = 12'b001101001100;
		14'b10010110101011: color_data = 12'b001101001100;
		14'b10010110101100: color_data = 12'b001101001100;
		14'b10010110101101: color_data = 12'b001101001100;
		14'b10010110101110: color_data = 12'b001101001100;
		14'b10010110101111: color_data = 12'b001101001100;
		14'b10010110110000: color_data = 12'b000000000000;
		14'b10011000010111: color_data = 12'b000000000000;
		14'b10011000011000: color_data = 12'b001101001100;
		14'b10011000011001: color_data = 12'b001101001100;
		14'b10011000011010: color_data = 12'b001101001100;
		14'b10011000011011: color_data = 12'b001101001100;
		14'b10011000011100: color_data = 12'b001101001100;
		14'b10011000011101: color_data = 12'b001101001100;
		14'b10011000011110: color_data = 12'b000000000000;
		14'b10011000101001: color_data = 12'b000000000000;
		14'b10011000101010: color_data = 12'b001101001100;
		14'b10011000101011: color_data = 12'b001101001100;
		14'b10011000101100: color_data = 12'b001101001100;
		14'b10011000101101: color_data = 12'b001101001100;
		14'b10011000101110: color_data = 12'b001101001100;
		14'b10011000101111: color_data = 12'b001101001100;
		14'b10011000110000: color_data = 12'b000000000000;
		14'b10011010010111: color_data = 12'b000000000000;
		14'b10011010011000: color_data = 12'b001101001100;
		14'b10011010011001: color_data = 12'b001101001100;
		14'b10011010011010: color_data = 12'b001101001100;
		14'b10011010011011: color_data = 12'b001101001100;
		14'b10011010011100: color_data = 12'b001101001100;
		14'b10011010011101: color_data = 12'b001101001100;
		14'b10011010011110: color_data = 12'b000000000000;
		14'b10011010101001: color_data = 12'b000000000000;
		14'b10011010101010: color_data = 12'b001101001100;
		14'b10011010101011: color_data = 12'b001101001100;
		14'b10011010101100: color_data = 12'b001101001100;
		14'b10011010101101: color_data = 12'b001101001100;
		14'b10011010101110: color_data = 12'b001101001100;
		14'b10011010101111: color_data = 12'b001101001100;
		14'b10011010110000: color_data = 12'b000000000000;
		14'b10011100010111: color_data = 12'b000000000000;
		14'b10011100011000: color_data = 12'b001101001100;
		14'b10011100011001: color_data = 12'b001101001100;
		14'b10011100011010: color_data = 12'b001101001100;
		14'b10011100011011: color_data = 12'b001101001100;
		14'b10011100011100: color_data = 12'b001101001100;
		14'b10011100011101: color_data = 12'b001101001100;
		14'b10011100011110: color_data = 12'b000000000000;
		14'b10011100101001: color_data = 12'b000000000000;
		14'b10011100101010: color_data = 12'b001101001100;
		14'b10011100101011: color_data = 12'b001101001100;
		14'b10011100101100: color_data = 12'b001101001100;
		14'b10011100101101: color_data = 12'b001101001100;
		14'b10011100101110: color_data = 12'b001101001100;
		14'b10011100101111: color_data = 12'b001101001100;
		14'b10011100110000: color_data = 12'b000000000000;
		14'b10011110010111: color_data = 12'b000000000000;
		14'b10011110011000: color_data = 12'b001101001100;
		14'b10011110011001: color_data = 12'b001101001100;
		14'b10011110011010: color_data = 12'b001101001100;
		14'b10011110011011: color_data = 12'b001101001100;
		14'b10011110011100: color_data = 12'b001101001100;
		14'b10011110011101: color_data = 12'b001101001100;
		14'b10011110011110: color_data = 12'b000000000000;
		14'b10011110101001: color_data = 12'b000000000000;
		14'b10011110101010: color_data = 12'b001101001100;
		14'b10011110101011: color_data = 12'b001101001100;
		14'b10011110101100: color_data = 12'b001101001100;
		14'b10011110101101: color_data = 12'b001101001100;
		14'b10011110101110: color_data = 12'b001101001100;
		14'b10011110101111: color_data = 12'b001101001100;
		14'b10011110110000: color_data = 12'b000000000000;
		14'b10100000010111: color_data = 12'b000000000000;
		14'b10100000011000: color_data = 12'b001101001100;
		14'b10100000011001: color_data = 12'b001101001100;
		14'b10100000011010: color_data = 12'b001101001100;
		14'b10100000011011: color_data = 12'b001101001100;
		14'b10100000011100: color_data = 12'b001101001100;
		14'b10100000011101: color_data = 12'b001101001100;
		14'b10100000011110: color_data = 12'b000000000000;
		14'b10100000101001: color_data = 12'b000000000000;
		14'b10100000101010: color_data = 12'b001101001100;
		14'b10100000101011: color_data = 12'b001101001100;
		14'b10100000101100: color_data = 12'b001101001100;
		14'b10100000101101: color_data = 12'b001101001100;
		14'b10100000101110: color_data = 12'b001101001100;
		14'b10100000101111: color_data = 12'b001101001100;
		14'b10100000110000: color_data = 12'b000000000000;
		14'b10100010010111: color_data = 12'b000000000000;
		14'b10100010011000: color_data = 12'b001101001100;
		14'b10100010011001: color_data = 12'b001101001100;
		14'b10100010011010: color_data = 12'b001101001100;
		14'b10100010011011: color_data = 12'b001101001100;
		14'b10100010011100: color_data = 12'b001101001100;
		14'b10100010011101: color_data = 12'b001101001100;
		14'b10100010011110: color_data = 12'b000000000000;
		14'b10100010101001: color_data = 12'b000000000000;
		14'b10100010101010: color_data = 12'b001101001100;
		14'b10100010101011: color_data = 12'b001101001100;
		14'b10100010101100: color_data = 12'b001101001100;
		14'b10100010101101: color_data = 12'b001101001100;
		14'b10100010101110: color_data = 12'b001101001100;
		14'b10100010101111: color_data = 12'b001101001100;
		14'b10100010110000: color_data = 12'b000000000000;
		14'b10100100010111: color_data = 12'b000000000000;
		14'b10100100011000: color_data = 12'b001101001100;
		14'b10100100011001: color_data = 12'b001101001100;
		14'b10100100011010: color_data = 12'b001101001100;
		14'b10100100011011: color_data = 12'b001101001100;
		14'b10100100011100: color_data = 12'b001101001100;
		14'b10100100011101: color_data = 12'b001101001100;
		14'b10100100011110: color_data = 12'b000000000000;
		14'b10100100101001: color_data = 12'b000000000000;
		14'b10100100101010: color_data = 12'b001101001100;
		14'b10100100101011: color_data = 12'b001101001100;
		14'b10100100101100: color_data = 12'b001101001100;
		14'b10100100101101: color_data = 12'b001101001100;
		14'b10100100101110: color_data = 12'b001101001100;
		14'b10100100101111: color_data = 12'b001101001100;
		14'b10100100110000: color_data = 12'b000000000000;
		14'b10100110001110: color_data = 12'b000000000000;
		14'b10100110001111: color_data = 12'b000000000000;
		14'b10100110010000: color_data = 12'b000000000000;
		14'b10100110010001: color_data = 12'b000000000000;
		14'b10100110010010: color_data = 12'b000000000000;
		14'b10100110010011: color_data = 12'b000000000000;
		14'b10100110010100: color_data = 12'b000000000000;
		14'b10100110010101: color_data = 12'b000000000000;
		14'b10100110010110: color_data = 12'b000000000000;
		14'b10100110010111: color_data = 12'b000000000000;
		14'b10100110011000: color_data = 12'b101101110101;
		14'b10100110011001: color_data = 12'b101101110101;
		14'b10100110011010: color_data = 12'b101101110101;
		14'b10100110011011: color_data = 12'b101101110101;
		14'b10100110011100: color_data = 12'b101101110101;
		14'b10100110011101: color_data = 12'b101101110101;
		14'b10100110011110: color_data = 12'b000000000000;
		14'b10100110101001: color_data = 12'b000000000000;
		14'b10100110101010: color_data = 12'b101101110101;
		14'b10100110101011: color_data = 12'b101101110101;
		14'b10100110101100: color_data = 12'b101101110101;
		14'b10100110101101: color_data = 12'b101101110101;
		14'b10100110101110: color_data = 12'b101101110101;
		14'b10100110101111: color_data = 12'b101101110101;
		14'b10100110110000: color_data = 12'b000000000000;
		14'b10100110110001: color_data = 12'b000000000000;
		14'b10100110110010: color_data = 12'b000000000000;
		14'b10100110110011: color_data = 12'b000000000000;
		14'b10100110110100: color_data = 12'b000000000000;
		14'b10100110110101: color_data = 12'b000000000000;
		14'b10100110110110: color_data = 12'b000000000000;
		14'b10100110110111: color_data = 12'b000000000000;
		14'b10100110111000: color_data = 12'b000000000000;
		14'b10100110111001: color_data = 12'b000000000000;
		14'b10100110111010: color_data = 12'b000000000000;
		14'b10100110111011: color_data = 12'b000000000000;
		14'b10101000001110: color_data = 12'b000000000000;
		14'b10101000001111: color_data = 12'b101101110101;
		14'b10101000010000: color_data = 12'b101101110101;
		14'b10101000010001: color_data = 12'b101101110101;
		14'b10101000010010: color_data = 12'b101101110101;
		14'b10101000010011: color_data = 12'b101101110101;
		14'b10101000010100: color_data = 12'b101101110101;
		14'b10101000010101: color_data = 12'b101101110101;
		14'b10101000010110: color_data = 12'b101101110101;
		14'b10101000010111: color_data = 12'b101101110101;
		14'b10101000011000: color_data = 12'b101101110101;
		14'b10101000011001: color_data = 12'b101101110101;
		14'b10101000011010: color_data = 12'b101101110101;
		14'b10101000011011: color_data = 12'b101101110101;
		14'b10101000011100: color_data = 12'b101101110101;
		14'b10101000011101: color_data = 12'b101101110101;
		14'b10101000011110: color_data = 12'b000000000000;
		14'b10101000101001: color_data = 12'b000000000000;
		14'b10101000101010: color_data = 12'b101101110101;
		14'b10101000101011: color_data = 12'b101101110101;
		14'b10101000101100: color_data = 12'b101101110101;
		14'b10101000101101: color_data = 12'b101101110101;
		14'b10101000101110: color_data = 12'b101101110101;
		14'b10101000101111: color_data = 12'b101101110101;
		14'b10101000110000: color_data = 12'b101101110101;
		14'b10101000110001: color_data = 12'b101101110101;
		14'b10101000110010: color_data = 12'b101101110101;
		14'b10101000110011: color_data = 12'b101101110101;
		14'b10101000110100: color_data = 12'b101101110101;
		14'b10101000110101: color_data = 12'b101101110101;
		14'b10101000110110: color_data = 12'b101101110101;
		14'b10101000110111: color_data = 12'b101101110101;
		14'b10101000111000: color_data = 12'b101101110101;
		14'b10101000111001: color_data = 12'b101101110101;
		14'b10101000111010: color_data = 12'b101101110101;
		14'b10101000111011: color_data = 12'b000000000000;
		14'b10101010001110: color_data = 12'b000000000000;
		14'b10101010001111: color_data = 12'b101101110101;
		14'b10101010010000: color_data = 12'b101101110101;
		14'b10101010010001: color_data = 12'b101101110101;
		14'b10101010010010: color_data = 12'b101101110101;
		14'b10101010010011: color_data = 12'b101101110101;
		14'b10101010010100: color_data = 12'b101101110101;
		14'b10101010010101: color_data = 12'b101101110101;
		14'b10101010010110: color_data = 12'b101101110101;
		14'b10101010010111: color_data = 12'b101101110101;
		14'b10101010011000: color_data = 12'b101101110101;
		14'b10101010011001: color_data = 12'b101101110101;
		14'b10101010011010: color_data = 12'b101101110101;
		14'b10101010011011: color_data = 12'b101101110101;
		14'b10101010011100: color_data = 12'b101101110101;
		14'b10101010011101: color_data = 12'b101101110101;
		14'b10101010011110: color_data = 12'b000000000000;
		14'b10101010101001: color_data = 12'b000000000000;
		14'b10101010101010: color_data = 12'b101101110101;
		14'b10101010101011: color_data = 12'b101101110101;
		14'b10101010101100: color_data = 12'b101101110101;
		14'b10101010101101: color_data = 12'b101101110101;
		14'b10101010101110: color_data = 12'b101101110101;
		14'b10101010101111: color_data = 12'b101101110101;
		14'b10101010110000: color_data = 12'b101101110101;
		14'b10101010110001: color_data = 12'b101101110101;
		14'b10101010110010: color_data = 12'b101101110101;
		14'b10101010110011: color_data = 12'b101101110101;
		14'b10101010110100: color_data = 12'b101101110101;
		14'b10101010110101: color_data = 12'b101101110101;
		14'b10101010110110: color_data = 12'b101101110101;
		14'b10101010110111: color_data = 12'b101101110101;
		14'b10101010111000: color_data = 12'b101101110101;
		14'b10101010111001: color_data = 12'b101101110101;
		14'b10101010111010: color_data = 12'b101101110101;
		14'b10101010111011: color_data = 12'b000000000000;
		14'b10101100001110: color_data = 12'b000000000000;
		14'b10101100001111: color_data = 12'b101101110101;
		14'b10101100010000: color_data = 12'b101101110101;
		14'b10101100010001: color_data = 12'b101101110101;
		14'b10101100010010: color_data = 12'b101101110101;
		14'b10101100010011: color_data = 12'b101101110101;
		14'b10101100010100: color_data = 12'b101101110101;
		14'b10101100010101: color_data = 12'b101101110101;
		14'b10101100010110: color_data = 12'b101101110101;
		14'b10101100010111: color_data = 12'b101101110101;
		14'b10101100011000: color_data = 12'b101101110101;
		14'b10101100011001: color_data = 12'b101101110101;
		14'b10101100011010: color_data = 12'b101101110101;
		14'b10101100011011: color_data = 12'b101101110101;
		14'b10101100011100: color_data = 12'b101101110101;
		14'b10101100011101: color_data = 12'b101101110101;
		14'b10101100011110: color_data = 12'b000000000000;
		14'b10101100101001: color_data = 12'b000000000000;
		14'b10101100101010: color_data = 12'b101101110101;
		14'b10101100101011: color_data = 12'b101101110101;
		14'b10101100101100: color_data = 12'b101101110101;
		14'b10101100101101: color_data = 12'b101101110101;
		14'b10101100101110: color_data = 12'b101101110101;
		14'b10101100101111: color_data = 12'b101101110101;
		14'b10101100110000: color_data = 12'b101101110101;
		14'b10101100110001: color_data = 12'b101101110101;
		14'b10101100110010: color_data = 12'b101101110101;
		14'b10101100110011: color_data = 12'b101101110101;
		14'b10101100110100: color_data = 12'b101101110101;
		14'b10101100110101: color_data = 12'b101101110101;
		14'b10101100110110: color_data = 12'b101101110101;
		14'b10101100110111: color_data = 12'b101101110101;
		14'b10101100111000: color_data = 12'b101101110101;
		14'b10101100111001: color_data = 12'b101101110101;
		14'b10101100111010: color_data = 12'b101101110101;
		14'b10101100111011: color_data = 12'b000000000000;
		14'b10101110001110: color_data = 12'b000000000000;
		14'b10101110001111: color_data = 12'b101101110101;
		14'b10101110010000: color_data = 12'b101101110101;
		14'b10101110010001: color_data = 12'b101101110101;
		14'b10101110010010: color_data = 12'b101101110101;
		14'b10101110010011: color_data = 12'b101101110101;
		14'b10101110010100: color_data = 12'b101101110101;
		14'b10101110010101: color_data = 12'b101101110101;
		14'b10101110010110: color_data = 12'b101101110101;
		14'b10101110010111: color_data = 12'b101101110101;
		14'b10101110011000: color_data = 12'b101101110101;
		14'b10101110011001: color_data = 12'b101101110101;
		14'b10101110011010: color_data = 12'b101101110101;
		14'b10101110011011: color_data = 12'b101101110101;
		14'b10101110011100: color_data = 12'b101101110101;
		14'b10101110011101: color_data = 12'b101101110101;
		14'b10101110011110: color_data = 12'b000000000000;
		14'b10101110101001: color_data = 12'b000000000000;
		14'b10101110101010: color_data = 12'b101101110101;
		14'b10101110101011: color_data = 12'b101101110101;
		14'b10101110101100: color_data = 12'b101101110101;
		14'b10101110101101: color_data = 12'b101101110101;
		14'b10101110101110: color_data = 12'b101101110101;
		14'b10101110101111: color_data = 12'b101101110101;
		14'b10101110110000: color_data = 12'b101101110101;
		14'b10101110110001: color_data = 12'b101101110101;
		14'b10101110110010: color_data = 12'b101101110101;
		14'b10101110110011: color_data = 12'b101101110101;
		14'b10101110110100: color_data = 12'b101101110101;
		14'b10101110110101: color_data = 12'b101101110101;
		14'b10101110110110: color_data = 12'b101101110101;
		14'b10101110110111: color_data = 12'b101101110101;
		14'b10101110111000: color_data = 12'b101101110101;
		14'b10101110111001: color_data = 12'b101101110101;
		14'b10101110111010: color_data = 12'b101101110101;
		14'b10101110111011: color_data = 12'b000000000000;
		14'b10110000001110: color_data = 12'b000000000000;
		14'b10110000001111: color_data = 12'b101101110101;
		14'b10110000010000: color_data = 12'b101101110101;
		14'b10110000010001: color_data = 12'b101101110101;
		14'b10110000010010: color_data = 12'b101101110101;
		14'b10110000010011: color_data = 12'b101101110101;
		14'b10110000010100: color_data = 12'b101101110101;
		14'b10110000010101: color_data = 12'b101101110101;
		14'b10110000010110: color_data = 12'b101101110101;
		14'b10110000010111: color_data = 12'b101101110101;
		14'b10110000011000: color_data = 12'b101101110101;
		14'b10110000011001: color_data = 12'b101101110101;
		14'b10110000011010: color_data = 12'b101101110101;
		14'b10110000011011: color_data = 12'b101101110101;
		14'b10110000011100: color_data = 12'b101101110101;
		14'b10110000011101: color_data = 12'b101101110101;
		14'b10110000011110: color_data = 12'b000000000000;
		14'b10110000101001: color_data = 12'b000000000000;
		14'b10110000101010: color_data = 12'b101101110101;
		14'b10110000101011: color_data = 12'b101101110101;
		14'b10110000101100: color_data = 12'b101101110101;
		14'b10110000101101: color_data = 12'b101101110101;
		14'b10110000101110: color_data = 12'b101101110101;
		14'b10110000101111: color_data = 12'b101101110101;
		14'b10110000110000: color_data = 12'b101101110101;
		14'b10110000110001: color_data = 12'b101101110101;
		14'b10110000110010: color_data = 12'b101101110101;
		14'b10110000110011: color_data = 12'b101101110101;
		14'b10110000110100: color_data = 12'b101101110101;
		14'b10110000110101: color_data = 12'b101101110101;
		14'b10110000110110: color_data = 12'b101101110101;
		14'b10110000110111: color_data = 12'b101101110101;
		14'b10110000111000: color_data = 12'b101101110101;
		14'b10110000111001: color_data = 12'b101101110101;
		14'b10110000111010: color_data = 12'b101101110101;
		14'b10110000111011: color_data = 12'b000000000000;
		14'b10110010001110: color_data = 12'b000000000000;
		14'b10110010001111: color_data = 12'b101101110101;
		14'b10110010010000: color_data = 12'b101101110101;
		14'b10110010010001: color_data = 12'b101101110101;
		14'b10110010010010: color_data = 12'b101101110101;
		14'b10110010010011: color_data = 12'b101101110101;
		14'b10110010010100: color_data = 12'b101101110101;
		14'b10110010010101: color_data = 12'b101101110101;
		14'b10110010010110: color_data = 12'b101101110101;
		14'b10110010010111: color_data = 12'b101101110101;
		14'b10110010011000: color_data = 12'b101101110101;
		14'b10110010011001: color_data = 12'b101101110101;
		14'b10110010011010: color_data = 12'b101101110101;
		14'b10110010011011: color_data = 12'b101101110101;
		14'b10110010011100: color_data = 12'b101101110101;
		14'b10110010011101: color_data = 12'b101101110101;
		14'b10110010011110: color_data = 12'b000000000000;
		14'b10110010101001: color_data = 12'b000000000000;
		14'b10110010101010: color_data = 12'b101101110101;
		14'b10110010101011: color_data = 12'b101101110101;
		14'b10110010101100: color_data = 12'b101101110101;
		14'b10110010101101: color_data = 12'b101101110101;
		14'b10110010101110: color_data = 12'b101101110101;
		14'b10110010101111: color_data = 12'b101101110101;
		14'b10110010110000: color_data = 12'b101101110101;
		14'b10110010110001: color_data = 12'b101101110101;
		14'b10110010110010: color_data = 12'b101101110101;
		14'b10110010110011: color_data = 12'b101101110101;
		14'b10110010110100: color_data = 12'b101101110101;
		14'b10110010110101: color_data = 12'b101101110101;
		14'b10110010110110: color_data = 12'b101101110101;
		14'b10110010110111: color_data = 12'b101101110101;
		14'b10110010111000: color_data = 12'b101101110101;
		14'b10110010111001: color_data = 12'b101101110101;
		14'b10110010111010: color_data = 12'b101101110101;
		14'b10110010111011: color_data = 12'b000000000000;
		14'b10110100001110: color_data = 12'b000000000000;
		14'b10110100001111: color_data = 12'b000000000000;
		14'b10110100010000: color_data = 12'b000000000000;
		14'b10110100010001: color_data = 12'b000000000000;
		14'b10110100010010: color_data = 12'b000000000000;
		14'b10110100010011: color_data = 12'b000000000000;
		14'b10110100010100: color_data = 12'b000000000000;
		14'b10110100010101: color_data = 12'b000000000000;
		14'b10110100010110: color_data = 12'b000000000000;
		14'b10110100010111: color_data = 12'b000000000000;
		14'b10110100011000: color_data = 12'b000000000000;
		14'b10110100011001: color_data = 12'b000000000000;
		14'b10110100011010: color_data = 12'b000000000000;
		14'b10110100011011: color_data = 12'b000000000000;
		14'b10110100011100: color_data = 12'b000000000000;
		14'b10110100011101: color_data = 12'b000000000000;
		14'b10110100011110: color_data = 12'b000000000000;
		14'b10110100101001: color_data = 12'b000000000000;
		14'b10110100101010: color_data = 12'b000000000000;
		14'b10110100101011: color_data = 12'b000000000000;
		14'b10110100101100: color_data = 12'b000000000000;
		14'b10110100101101: color_data = 12'b000000000000;
		14'b10110100101110: color_data = 12'b000000000000;
		14'b10110100101111: color_data = 12'b000000000000;
		14'b10110100110000: color_data = 12'b000000000000;
		14'b10110100110001: color_data = 12'b000000000000;
		14'b10110100110010: color_data = 12'b000000000000;
		14'b10110100110011: color_data = 12'b000000000000;
		14'b10110100110100: color_data = 12'b000000000000;
		14'b10110100110101: color_data = 12'b000000000000;
		14'b10110100110110: color_data = 12'b000000000000;
		14'b10110100110111: color_data = 12'b000000000000;
		14'b10110100111000: color_data = 12'b000000000000;
		14'b10110100111001: color_data = 12'b000000000000;
		14'b10110100111010: color_data = 12'b000000000000;
		14'b10110100111011: color_data = 12'b000000000000;
        default: color_data = 12'b111111111111;
	endcase
endmodule