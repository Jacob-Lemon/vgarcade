`timescale 1ns / 1ps
module orange_rom (
    input wire clk,
    input wire [5:0] row,
    input wire [5:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 40 + col) >= 0 && (row * 40 + col) <= 60) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 61 && (row * 40 + col) <= 71) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 72 && (row * 40 + col) <= 97) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 98 && (row * 40 + col) <= 100) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 101 && (row * 40 + col) <= 111) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 112 && (row * 40 + col) <= 114) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 115 && (row * 40 + col) <= 134) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 135 && (row * 40 + col) <= 137) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 138 && (row * 40 + col) <= 154) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 155 && (row * 40 + col) <= 156) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 157 && (row * 40 + col) <= 173) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 174 && (row * 40 + col) <= 175) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 176 && (row * 40 + col) <= 196) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 197 && (row * 40 + col) <= 197) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 198 && (row * 40 + col) <= 213) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 214 && (row * 40 + col) <= 214) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 215 && (row * 40 + col) <= 237) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 238 && (row * 40 + col) <= 238) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 239 && (row * 40 + col) <= 253) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 254 && (row * 40 + col) <= 254) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 255 && (row * 40 + col) <= 277) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 278 && (row * 40 + col) <= 278) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 279 && (row * 40 + col) <= 293) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 294 && (row * 40 + col) <= 295) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 296 && (row * 40 + col) <= 316) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 317 && (row * 40 + col) <= 317) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 318 && (row * 40 + col) <= 333) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 334 && (row * 40 + col) <= 334) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 335 && (row * 40 + col) <= 335) color_data <= 12'b101101110101; else
        if ((row * 40 + col) >= 336 && (row * 40 + col) <= 337) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 338 && (row * 40 + col) <= 354) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 355 && (row * 40 + col) <= 356) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 357 && (row * 40 + col) <= 371) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 372 && (row * 40 + col) <= 374) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 375 && (row * 40 + col) <= 375) color_data <= 12'b101101110101; else
        if ((row * 40 + col) >= 376 && (row * 40 + col) <= 380) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 381 && (row * 40 + col) <= 391) color_data <= 12'b001010110000; else
        if ((row * 40 + col) >= 392 && (row * 40 + col) <= 394) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 395 && (row * 40 + col) <= 408) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 409 && (row * 40 + col) <= 411) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 412 && (row * 40 + col) <= 413) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 414 && (row * 40 + col) <= 414) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 415 && (row * 40 + col) <= 415) color_data <= 12'b101101110101; else
        if ((row * 40 + col) >= 416 && (row * 40 + col) <= 416) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 417 && (row * 40 + col) <= 418) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 419 && (row * 40 + col) <= 431) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 432 && (row * 40 + col) <= 446) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 447 && (row * 40 + col) <= 448) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 449 && (row * 40 + col) <= 453) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 454 && (row * 40 + col) <= 454) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 455 && (row * 40 + col) <= 455) color_data <= 12'b101101110101; else
        if ((row * 40 + col) >= 456 && (row * 40 + col) <= 456) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 457 && (row * 40 + col) <= 461) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 462 && (row * 40 + col) <= 463) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 464 && (row * 40 + col) <= 485) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 486 && (row * 40 + col) <= 486) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 487 && (row * 40 + col) <= 493) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 494 && (row * 40 + col) <= 494) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 495 && (row * 40 + col) <= 495) color_data <= 12'b101101110101; else
        if ((row * 40 + col) >= 496 && (row * 40 + col) <= 496) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 497 && (row * 40 + col) <= 503) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 504 && (row * 40 + col) <= 504) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 505 && (row * 40 + col) <= 524) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 525 && (row * 40 + col) <= 525) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 526 && (row * 40 + col) <= 533) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 534 && (row * 40 + col) <= 535) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 536 && (row * 40 + col) <= 544) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 545 && (row * 40 + col) <= 545) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 546 && (row * 40 + col) <= 563) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 564 && (row * 40 + col) <= 564) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 565 && (row * 40 + col) <= 574) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 575 && (row * 40 + col) <= 575) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 576 && (row * 40 + col) <= 585) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 586 && (row * 40 + col) <= 586) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 587 && (row * 40 + col) <= 602) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 603 && (row * 40 + col) <= 603) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 604 && (row * 40 + col) <= 626) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 627 && (row * 40 + col) <= 627) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 628 && (row * 40 + col) <= 641) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 642 && (row * 40 + col) <= 642) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 643 && (row * 40 + col) <= 667) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 668 && (row * 40 + col) <= 668) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 669 && (row * 40 + col) <= 681) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 682 && (row * 40 + col) <= 682) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 683 && (row * 40 + col) <= 707) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 708 && (row * 40 + col) <= 708) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 709 && (row * 40 + col) <= 720) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 721 && (row * 40 + col) <= 721) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 722 && (row * 40 + col) <= 748) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 749 && (row * 40 + col) <= 749) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 750 && (row * 40 + col) <= 760) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 761 && (row * 40 + col) <= 761) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 762 && (row * 40 + col) <= 788) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 789 && (row * 40 + col) <= 789) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 790 && (row * 40 + col) <= 800) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 801 && (row * 40 + col) <= 801) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 802 && (row * 40 + col) <= 828) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 829 && (row * 40 + col) <= 829) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 830 && (row * 40 + col) <= 839) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 840 && (row * 40 + col) <= 840) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 841 && (row * 40 + col) <= 869) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 870 && (row * 40 + col) <= 870) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 871 && (row * 40 + col) <= 879) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 880 && (row * 40 + col) <= 880) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 881 && (row * 40 + col) <= 909) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 910 && (row * 40 + col) <= 910) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 911 && (row * 40 + col) <= 919) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 920 && (row * 40 + col) <= 920) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 921 && (row * 40 + col) <= 949) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 950 && (row * 40 + col) <= 950) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 951 && (row * 40 + col) <= 959) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 960 && (row * 40 + col) <= 960) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 961 && (row * 40 + col) <= 989) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 990 && (row * 40 + col) <= 990) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 991 && (row * 40 + col) <= 999) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1000 && (row * 40 + col) <= 1000) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1001 && (row * 40 + col) <= 1029) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1030 && (row * 40 + col) <= 1030) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1031 && (row * 40 + col) <= 1039) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1040 && (row * 40 + col) <= 1040) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1041 && (row * 40 + col) <= 1069) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1070 && (row * 40 + col) <= 1070) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1071 && (row * 40 + col) <= 1079) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1080 && (row * 40 + col) <= 1080) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1081 && (row * 40 + col) <= 1109) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1110 && (row * 40 + col) <= 1110) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1111 && (row * 40 + col) <= 1120) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1121 && (row * 40 + col) <= 1121) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1122 && (row * 40 + col) <= 1148) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1149 && (row * 40 + col) <= 1149) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1150 && (row * 40 + col) <= 1160) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1161 && (row * 40 + col) <= 1161) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1162 && (row * 40 + col) <= 1188) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1189 && (row * 40 + col) <= 1189) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1190 && (row * 40 + col) <= 1200) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1201 && (row * 40 + col) <= 1201) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1202 && (row * 40 + col) <= 1228) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1229 && (row * 40 + col) <= 1229) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1230 && (row * 40 + col) <= 1241) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1242 && (row * 40 + col) <= 1242) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1243 && (row * 40 + col) <= 1267) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1268 && (row * 40 + col) <= 1268) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1269 && (row * 40 + col) <= 1281) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1282 && (row * 40 + col) <= 1282) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1283 && (row * 40 + col) <= 1307) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1308 && (row * 40 + col) <= 1308) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1309 && (row * 40 + col) <= 1322) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1323 && (row * 40 + col) <= 1323) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1324 && (row * 40 + col) <= 1346) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1347 && (row * 40 + col) <= 1347) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1348 && (row * 40 + col) <= 1363) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1364 && (row * 40 + col) <= 1364) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1365 && (row * 40 + col) <= 1385) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1386 && (row * 40 + col) <= 1386) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1387 && (row * 40 + col) <= 1404) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1405 && (row * 40 + col) <= 1405) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1406 && (row * 40 + col) <= 1424) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1425 && (row * 40 + col) <= 1425) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1426 && (row * 40 + col) <= 1445) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1446 && (row * 40 + col) <= 1446) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1447 && (row * 40 + col) <= 1463) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1464 && (row * 40 + col) <= 1464) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1465 && (row * 40 + col) <= 1486) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1487 && (row * 40 + col) <= 1488) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1489 && (row * 40 + col) <= 1501) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1502 && (row * 40 + col) <= 1503) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1504 && (row * 40 + col) <= 1528) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1529 && (row * 40 + col) <= 1531) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1532 && (row * 40 + col) <= 1538) color_data <= 12'b111110110000; else
        if ((row * 40 + col) >= 1539 && (row * 40 + col) <= 1541) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1542 && (row * 40 + col) <= 1571) color_data <= 12'b111111111111; else
        if ((row * 40 + col) >= 1572 && (row * 40 + col) <= 1578) color_data <= 12'b000000000000; else
        if ((row * 40 + col) >= 1579 && (row * 40 + col) < 1600) color_data <= 12'b111111111111; else
        color_data <= 12'b000000000000;
    end
endmodule
