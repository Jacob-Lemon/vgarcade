module joystick_rom (
    input wire clk,
    input wire [6:0] row,
    input wire [6:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 70 + col) >= 0 && (row * 70 + col) <= 96) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 97 && (row * 70 + col) <= 112) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 113 && (row * 70 + col) <= 163) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 164 && (row * 70 + col) <= 185) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 186 && (row * 70 + col) <= 230) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 231 && (row * 70 + col) <= 258) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 259 && (row * 70 + col) <= 298) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 299 && (row * 70 + col) <= 330) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 331 && (row * 70 + col) <= 366) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 367 && (row * 70 + col) <= 402) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 403 && (row * 70 + col) <= 435) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 436 && (row * 70 + col) <= 473) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 474 && (row * 70 + col) <= 503) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 504 && (row * 70 + col) <= 545) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 546 && (row * 70 + col) <= 572) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 573 && (row * 70 + col) <= 616) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 617 && (row * 70 + col) <= 641) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 642 && (row * 70 + col) <= 657) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 658 && (row * 70 + col) <= 671) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 672 && (row * 70 + col) <= 687) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 688 && (row * 70 + col) <= 710) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 711 && (row * 70 + col) <= 724) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 725 && (row * 70 + col) <= 744) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 745 && (row * 70 + col) <= 758) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 759 && (row * 70 + col) <= 779) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 780 && (row * 70 + col) <= 792) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 793 && (row * 70 + col) <= 816) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 817 && (row * 70 + col) <= 829) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 830 && (row * 70 + col) <= 848) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 849 && (row * 70 + col) <= 860) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 861 && (row * 70 + col) <= 888) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 889 && (row * 70 + col) <= 900) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 901 && (row * 70 + col) <= 917) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 918 && (row * 70 + col) <= 929) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 930 && (row * 70 + col) <= 959) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 960 && (row * 70 + col) <= 971) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 972 && (row * 70 + col) <= 986) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 987 && (row * 70 + col) <= 997) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 998 && (row * 70 + col) <= 1031) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1032 && (row * 70 + col) <= 1042) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1043 && (row * 70 + col) <= 1056) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1057 && (row * 70 + col) <= 1066) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1067 && (row * 70 + col) <= 1102) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1103 && (row * 70 + col) <= 1113) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1114 && (row * 70 + col) <= 1125) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1126 && (row * 70 + col) <= 1135) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1136 && (row * 70 + col) <= 1173) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1174 && (row * 70 + col) <= 1183) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1184 && (row * 70 + col) <= 1194) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1195 && (row * 70 + col) <= 1204) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1205 && (row * 70 + col) <= 1244) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1245 && (row * 70 + col) <= 1254) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1255 && (row * 70 + col) <= 1264) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1265 && (row * 70 + col) <= 1273) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1274 && (row * 70 + col) <= 1315) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1316 && (row * 70 + col) <= 1324) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1325 && (row * 70 + col) <= 1333) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1334 && (row * 70 + col) <= 1343) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1344 && (row * 70 + col) <= 1385) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1386 && (row * 70 + col) <= 1395) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1396 && (row * 70 + col) <= 1403) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1404 && (row * 70 + col) <= 1412) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1413 && (row * 70 + col) <= 1456) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1457 && (row * 70 + col) <= 1465) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1466 && (row * 70 + col) <= 1472) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1473 && (row * 70 + col) <= 1481) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1482 && (row * 70 + col) <= 1527) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1528 && (row * 70 + col) <= 1536) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1537 && (row * 70 + col) <= 1542) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1543 && (row * 70 + col) <= 1551) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1552 && (row * 70 + col) <= 1597) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1598 && (row * 70 + col) <= 1606) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1607 && (row * 70 + col) <= 1612) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1613 && (row * 70 + col) <= 1620) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1621 && (row * 70 + col) <= 1668) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1669 && (row * 70 + col) <= 1676) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1677 && (row * 70 + col) <= 1681) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1682 && (row * 70 + col) <= 1690) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1691 && (row * 70 + col) <= 1738) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1739 && (row * 70 + col) <= 1747) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1748 && (row * 70 + col) <= 1751) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1752 && (row * 70 + col) <= 1759) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1760 && (row * 70 + col) <= 1809) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1810 && (row * 70 + col) <= 1817) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1818 && (row * 70 + col) <= 1821) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1822 && (row * 70 + col) <= 1829) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1830 && (row * 70 + col) <= 1879) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1880 && (row * 70 + col) <= 1887) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1888 && (row * 70 + col) <= 1890) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1891 && (row * 70 + col) <= 1899) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1900 && (row * 70 + col) <= 1949) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 1950 && (row * 70 + col) <= 1958) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1959 && (row * 70 + col) <= 1960) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 1961 && (row * 70 + col) <= 1968) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 1969 && (row * 70 + col) <= 2020) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2021 && (row * 70 + col) <= 2028) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2029 && (row * 70 + col) <= 2030) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2031 && (row * 70 + col) <= 2038) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2039 && (row * 70 + col) <= 2090) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2091 && (row * 70 + col) <= 2098) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2099 && (row * 70 + col) <= 2100) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2101 && (row * 70 + col) <= 2108) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2109 && (row * 70 + col) <= 2160) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2161 && (row * 70 + col) <= 2168) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2169 && (row * 70 + col) <= 2170) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2171 && (row * 70 + col) <= 2178) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2179 && (row * 70 + col) <= 2230) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2231 && (row * 70 + col) <= 2238) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2239 && (row * 70 + col) <= 2240) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2241 && (row * 70 + col) <= 2248) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2249 && (row * 70 + col) <= 2300) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2301 && (row * 70 + col) <= 2308) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2309 && (row * 70 + col) <= 2310) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2311 && (row * 70 + col) <= 2318) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2319 && (row * 70 + col) <= 2370) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2371 && (row * 70 + col) <= 2378) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2379 && (row * 70 + col) <= 2380) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2381 && (row * 70 + col) <= 2388) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2389 && (row * 70 + col) <= 2440) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2441 && (row * 70 + col) <= 2448) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2449 && (row * 70 + col) <= 2450) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2451 && (row * 70 + col) <= 2458) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2459 && (row * 70 + col) <= 2510) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2511 && (row * 70 + col) <= 2518) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2519 && (row * 70 + col) <= 2520) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2521 && (row * 70 + col) <= 2528) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2529 && (row * 70 + col) <= 2580) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2581 && (row * 70 + col) <= 2588) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2589 && (row * 70 + col) <= 2590) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2591 && (row * 70 + col) <= 2598) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2599 && (row * 70 + col) <= 2650) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2651 && (row * 70 + col) <= 2658) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2659 && (row * 70 + col) <= 2660) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2661 && (row * 70 + col) <= 2668) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2669 && (row * 70 + col) <= 2720) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2721 && (row * 70 + col) <= 2728) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2729 && (row * 70 + col) <= 2730) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2731 && (row * 70 + col) <= 2738) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2739 && (row * 70 + col) <= 2790) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2791 && (row * 70 + col) <= 2798) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2799 && (row * 70 + col) <= 2800) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2801 && (row * 70 + col) <= 2808) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2809 && (row * 70 + col) <= 2860) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2861 && (row * 70 + col) <= 2868) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2869 && (row * 70 + col) <= 2870) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2871 && (row * 70 + col) <= 2878) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2879 && (row * 70 + col) <= 2930) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 2931 && (row * 70 + col) <= 2938) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2939 && (row * 70 + col) <= 2940) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 2941 && (row * 70 + col) <= 2949) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 2950 && (row * 70 + col) <= 2999) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3000 && (row * 70 + col) <= 3008) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3009 && (row * 70 + col) <= 3011) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3012 && (row * 70 + col) <= 3019) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3020 && (row * 70 + col) <= 3069) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3070 && (row * 70 + col) <= 3077) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3078 && (row * 70 + col) <= 3081) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3082 && (row * 70 + col) <= 3089) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3090 && (row * 70 + col) <= 3139) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3140 && (row * 70 + col) <= 3147) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3148 && (row * 70 + col) <= 3151) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3152 && (row * 70 + col) <= 3160) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3161 && (row * 70 + col) <= 3208) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3209 && (row * 70 + col) <= 3217) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3218 && (row * 70 + col) <= 3222) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3223 && (row * 70 + col) <= 3230) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3231 && (row * 70 + col) <= 3278) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3279 && (row * 70 + col) <= 3286) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3287 && (row * 70 + col) <= 3292) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3293 && (row * 70 + col) <= 3301) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3302 && (row * 70 + col) <= 3347) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3348 && (row * 70 + col) <= 3356) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3357 && (row * 70 + col) <= 3362) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3363 && (row * 70 + col) <= 3371) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3372 && (row * 70 + col) <= 3417) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3418 && (row * 70 + col) <= 3426) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3427 && (row * 70 + col) <= 3433) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3434 && (row * 70 + col) <= 3442) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3443 && (row * 70 + col) <= 3486) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3487 && (row * 70 + col) <= 3495) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3496 && (row * 70 + col) <= 3503) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3504 && (row * 70 + col) <= 3513) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3514 && (row * 70 + col) <= 3555) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3556 && (row * 70 + col) <= 3565) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3566 && (row * 70 + col) <= 3574) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3575 && (row * 70 + col) <= 3583) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3584 && (row * 70 + col) <= 3625) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3626 && (row * 70 + col) <= 3634) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3635 && (row * 70 + col) <= 3644) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3645 && (row * 70 + col) <= 3654) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3655 && (row * 70 + col) <= 3694) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3695 && (row * 70 + col) <= 3704) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3705 && (row * 70 + col) <= 3715) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3716 && (row * 70 + col) <= 3725) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3726 && (row * 70 + col) <= 3763) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3764 && (row * 70 + col) <= 3773) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3774 && (row * 70 + col) <= 3786) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3787 && (row * 70 + col) <= 3796) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3797 && (row * 70 + col) <= 3832) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3833 && (row * 70 + col) <= 3843) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3844 && (row * 70 + col) <= 3856) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3857 && (row * 70 + col) <= 3867) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3868 && (row * 70 + col) <= 3901) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3902 && (row * 70 + col) <= 3912) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3913 && (row * 70 + col) <= 3927) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3928 && (row * 70 + col) <= 3939) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3940 && (row * 70 + col) <= 3969) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 3970 && (row * 70 + col) <= 3981) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 3982 && (row * 70 + col) <= 3998) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 3999 && (row * 70 + col) <= 4010) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4011 && (row * 70 + col) <= 4038) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 4039 && (row * 70 + col) <= 4050) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4051 && (row * 70 + col) <= 4069) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4070 && (row * 70 + col) <= 4082) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4083 && (row * 70 + col) <= 4106) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 4107 && (row * 70 + col) <= 4119) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4120 && (row * 70 + col) <= 4140) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4141 && (row * 70 + col) <= 4154) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4155 && (row * 70 + col) <= 4174) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 4175 && (row * 70 + col) <= 4188) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4189 && (row * 70 + col) <= 4211) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4212 && (row * 70 + col) <= 4227) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4228 && (row * 70 + col) <= 4241) color_data <= 12'b100010001000; else
        if ((row * 70 + col) >= 4242 && (row * 70 + col) <= 4257) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4258 && (row * 70 + col) <= 4282) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4283 && (row * 70 + col) <= 4326) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4327 && (row * 70 + col) <= 4353) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4354 && (row * 70 + col) <= 4395) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4396 && (row * 70 + col) <= 4424) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4425 && (row * 70 + col) <= 4464) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4465 && (row * 70 + col) <= 4496) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4497 && (row * 70 + col) <= 4532) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4533 && (row * 70 + col) <= 4568) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4569 && (row * 70 + col) <= 4600) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4601 && (row * 70 + col) <= 4640) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4641 && (row * 70 + col) <= 4668) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4669 && (row * 70 + col) <= 4713) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4714 && (row * 70 + col) <= 4735) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4736 && (row * 70 + col) <= 4786) color_data <= 12'b000000000000; else
        if ((row * 70 + col) >= 4787 && (row * 70 + col) <= 4802) color_data <= 12'b111111111111; else
        if ((row * 70 + col) >= 4803 && (row * 70 + col) < 4900) color_data <= 12'b000000000000; else
        color_data <= 12'b000000000000;
    end
endmodule
