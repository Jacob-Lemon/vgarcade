`timescale 1ns / 1ps
module killscreen_rom (
    input wire clk,
    input wire [8:0] row,
    input wire [9:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 640 + col) >= 0 && (row * 640 + col) <= 8518) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 8519 && (row * 640 + col) <= 8533) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 8534 && (row * 640 + col) <= 9156) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 9157 && (row * 640 + col) <= 9175) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 9176 && (row * 640 + col) <= 9794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 9795 && (row * 640 + col) <= 9817) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 9818 && (row * 640 + col) <= 10431) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 10432 && (row * 640 + col) <= 10460) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 10461 && (row * 640 + col) <= 11071) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 11072 && (row * 640 + col) <= 11100) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 11101 && (row * 640 + col) <= 11710) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 11711 && (row * 640 + col) <= 11741) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 11742 && (row * 640 + col) <= 12348) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 12349 && (row * 640 + col) <= 12383) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 12384 && (row * 640 + col) <= 12988) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 12989 && (row * 640 + col) <= 13023) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 13024 && (row * 640 + col) <= 13627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 13628 && (row * 640 + col) <= 13664) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 13665 && (row * 640 + col) <= 14265) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 14266 && (row * 640 + col) <= 14306) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 14307 && (row * 640 + col) <= 14905) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 14906 && (row * 640 + col) <= 14946) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 14947 && (row * 640 + col) <= 15545) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 15546 && (row * 640 + col) <= 15586) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 15587 && (row * 640 + col) <= 16184) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 16185 && (row * 640 + col) <= 16227) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 16228 && (row * 640 + col) <= 16824) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 16825 && (row * 640 + col) <= 16867) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 16868 && (row * 640 + col) <= 17463) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 17464 && (row * 640 + col) <= 17508) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 17509 && (row * 640 + col) <= 18103) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 18104 && (row * 640 + col) <= 18148) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 18149 && (row * 640 + col) <= 18742) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 18743 && (row * 640 + col) <= 18789) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 18790 && (row * 640 + col) <= 19382) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 19383 && (row * 640 + col) <= 19429) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 19430 && (row * 640 + col) <= 20022) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 20023 && (row * 640 + col) <= 20069) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 20070 && (row * 640 + col) <= 20662) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 20663 && (row * 640 + col) <= 20709) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 20710 && (row * 640 + col) <= 21302) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 21303 && (row * 640 + col) <= 21349) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 21350 && (row * 640 + col) <= 21942) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 21943 && (row * 640 + col) <= 21989) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 21990 && (row * 640 + col) <= 22582) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 22583 && (row * 640 + col) <= 22629) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 22630 && (row * 640 + col) <= 23222) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 23223 && (row * 640 + col) <= 23269) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 23270 && (row * 640 + col) <= 23862) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 23863 && (row * 640 + col) <= 23909) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 23910 && (row * 640 + col) <= 24502) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 24503 && (row * 640 + col) <= 24549) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 24550 && (row * 640 + col) <= 25142) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 25143 && (row * 640 + col) <= 25189) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 25190 && (row * 640 + col) <= 25782) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 25783 && (row * 640 + col) <= 25829) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 25830 && (row * 640 + col) <= 26422) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 26423 && (row * 640 + col) <= 26469) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 26470 && (row * 640 + col) <= 27062) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 27063 && (row * 640 + col) <= 27109) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 27110 && (row * 640 + col) <= 27703) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 27704 && (row * 640 + col) <= 27749) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 27750 && (row * 640 + col) <= 28343) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 28344 && (row * 640 + col) <= 28388) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 28389 && (row * 640 + col) <= 28984) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 28985 && (row * 640 + col) <= 29028) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 29029 && (row * 640 + col) <= 29624) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 29625 && (row * 640 + col) <= 29667) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 29668 && (row * 640 + col) <= 30265) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 30266 && (row * 640 + col) <= 30307) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 30308 && (row * 640 + col) <= 30905) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 30906 && (row * 640 + col) <= 30946) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 30947 && (row * 640 + col) <= 31545) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 31546 && (row * 640 + col) <= 31586) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 31587 && (row * 640 + col) <= 32186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 32187 && (row * 640 + col) <= 32225) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 32226 && (row * 640 + col) <= 32828) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 32829 && (row * 640 + col) <= 32864) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 32865 && (row * 640 + col) <= 33468) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 33469 && (row * 640 + col) <= 33503) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 33504 && (row * 640 + col) <= 34109) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 34110 && (row * 640 + col) <= 34143) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 34144 && (row * 640 + col) <= 34751) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 34752 && (row * 640 + col) <= 34781) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 34782 && (row * 640 + col) <= 35391) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 35392 && (row * 640 + col) <= 35420) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 35421 && (row * 640 + col) <= 36032) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 36033 && (row * 640 + col) <= 36059) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 36060 && (row * 640 + col) <= 36674) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 36675 && (row * 640 + col) <= 36697) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 36698 && (row * 640 + col) <= 37316) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 37317 && (row * 640 + col) <= 37335) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 37336 && (row * 640 + col) <= 37958) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 37959 && (row * 640 + col) <= 37973) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 37974 && (row * 640 + col) <= 41998) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 41999 && (row * 640 + col) <= 42001) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 42002 && (row * 640 + col) <= 42638) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 42639 && (row * 640 + col) <= 42641) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 42642 && (row * 640 + col) <= 43278) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 43279 && (row * 640 + col) <= 43281) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 43282 && (row * 640 + col) <= 43918) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 43919 && (row * 640 + col) <= 43921) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 43922 && (row * 640 + col) <= 44558) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 44559 && (row * 640 + col) <= 44561) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 44562 && (row * 640 + col) <= 45198) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 45199 && (row * 640 + col) <= 45201) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 45202 && (row * 640 + col) <= 45439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 45440 && (row * 640 + col) <= 45445) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 45446 && (row * 640 + col) <= 45838) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 45839 && (row * 640 + col) <= 45841) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 45842 && (row * 640 + col) <= 46079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 46080 && (row * 640 + col) <= 46085) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46086 && (row * 640 + col) <= 46478) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 46479 && (row * 640 + col) <= 46481) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 46482 && (row * 640 + col) <= 46719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 46720 && (row * 640 + col) <= 46726) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 46727 && (row * 640 + col) <= 47118) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 47119 && (row * 640 + col) <= 47121) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 47122 && (row * 640 + col) <= 47359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 47360 && (row * 640 + col) <= 47379) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 47380 && (row * 640 + col) <= 47758) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 47759 && (row * 640 + col) <= 47761) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 47762 && (row * 640 + col) <= 47999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 48000 && (row * 640 + col) <= 48019) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48020 && (row * 640 + col) <= 48398) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 48399 && (row * 640 + col) <= 48401) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 48402 && (row * 640 + col) <= 48639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 48640 && (row * 640 + col) <= 48664) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 48665 && (row * 640 + col) <= 49038) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 49039 && (row * 640 + col) <= 49041) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 49042 && (row * 640 + col) <= 49279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 49280 && (row * 640 + col) <= 49305) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49306 && (row * 640 + col) <= 49678) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 49679 && (row * 640 + col) <= 49681) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 49682 && (row * 640 + col) <= 49919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 49920 && (row * 640 + col) <= 49945) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 49946 && (row * 640 + col) <= 50318) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 50319 && (row * 640 + col) <= 50321) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 50322 && (row * 640 + col) <= 50559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 50560 && (row * 640 + col) <= 50587) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 50588 && (row * 640 + col) <= 50958) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 50959 && (row * 640 + col) <= 50961) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 50962 && (row * 640 + col) <= 51199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 51200 && (row * 640 + col) <= 51230) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51231 && (row * 640 + col) <= 51598) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 51599 && (row * 640 + col) <= 51601) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 51602 && (row * 640 + col) <= 51839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 51840 && (row * 640 + col) <= 51871) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 51872 && (row * 640 + col) <= 52238) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 52239 && (row * 640 + col) <= 52241) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 52242 && (row * 640 + col) <= 52479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 52480 && (row * 640 + col) <= 52512) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 52513 && (row * 640 + col) <= 52878) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 52879 && (row * 640 + col) <= 52881) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 52882 && (row * 640 + col) <= 53119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 53120 && (row * 640 + col) <= 53153) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53154 && (row * 640 + col) <= 53518) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 53519 && (row * 640 + col) <= 53521) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 53522 && (row * 640 + col) <= 53759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 53760 && (row * 640 + col) <= 53794) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 53795 && (row * 640 + col) <= 54158) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 54159 && (row * 640 + col) <= 54161) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 54162 && (row * 640 + col) <= 54399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 54400 && (row * 640 + col) <= 54453) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 54454 && (row * 640 + col) <= 54798) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 54799 && (row * 640 + col) <= 54801) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 54802 && (row * 640 + col) <= 55039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 55040 && (row * 640 + col) <= 55093) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55094 && (row * 640 + col) <= 55438) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 55439 && (row * 640 + col) <= 55441) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 55442 && (row * 640 + col) <= 55679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 55680 && (row * 640 + col) <= 55734) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 55735 && (row * 640 + col) <= 56078) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 56079 && (row * 640 + col) <= 56081) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56082 && (row * 640 + col) <= 56319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 56320 && (row * 640 + col) <= 56379) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 56380 && (row * 640 + col) <= 56718) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 56719 && (row * 640 + col) <= 56721) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 56722 && (row * 640 + col) <= 56959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 56960 && (row * 640 + col) <= 57019) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57020 && (row * 640 + col) <= 57358) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 57359 && (row * 640 + col) <= 57361) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 57362 && (row * 640 + col) <= 57599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 57600 && (row * 640 + col) <= 57659) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 57660 && (row * 640 + col) <= 57998) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 57999 && (row * 640 + col) <= 58001) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58002 && (row * 640 + col) <= 58239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 58240 && (row * 640 + col) <= 58307) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58308 && (row * 640 + col) <= 58638) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 58639 && (row * 640 + col) <= 58641) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 58642 && (row * 640 + col) <= 58879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 58880 && (row * 640 + col) <= 58948) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 58949 && (row * 640 + col) <= 59278) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 59279 && (row * 640 + col) <= 59281) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59282 && (row * 640 + col) <= 59519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 59520 && (row * 640 + col) <= 59588) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 59589 && (row * 640 + col) <= 59918) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 59919 && (row * 640 + col) <= 59921) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 59922 && (row * 640 + col) <= 60159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 60160 && (row * 640 + col) <= 60239) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60240 && (row * 640 + col) <= 60558) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 60559 && (row * 640 + col) <= 60561) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 60562 && (row * 640 + col) <= 60799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 60800 && (row * 640 + col) <= 60879) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 60880 && (row * 640 + col) <= 61198) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 61199 && (row * 640 + col) <= 61201) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61202 && (row * 640 + col) <= 61439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 61440 && (row * 640 + col) <= 61518) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 61519 && (row * 640 + col) <= 61838) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 61839 && (row * 640 + col) <= 61841) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 61842 && (row * 640 + col) <= 62079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 62080 && (row * 640 + col) <= 62142) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62143 && (row * 640 + col) <= 62478) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 62479 && (row * 640 + col) <= 62481) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 62482 && (row * 640 + col) <= 62532) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 62533 && (row * 640 + col) <= 62547) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62548 && (row * 640 + col) <= 62719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 62720 && (row * 640 + col) <= 62782) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 62783 && (row * 640 + col) <= 63118) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 63119 && (row * 640 + col) <= 63121) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63122 && (row * 640 + col) <= 63172) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 63173 && (row * 640 + col) <= 63187) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63188 && (row * 640 + col) <= 63359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 63360 && (row * 640 + col) <= 63400) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63401 && (row * 640 + col) <= 63758) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 63759 && (row * 640 + col) <= 63761) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 63762 && (row * 640 + col) <= 63811) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 63812 && (row * 640 + col) <= 63837) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 63838 && (row * 640 + col) <= 63999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 64000 && (row * 640 + col) <= 64039) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64040 && (row * 640 + col) <= 64398) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 64399 && (row * 640 + col) <= 64401) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 64402 && (row * 640 + col) <= 64450) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 64451 && (row * 640 + col) <= 64478) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64479 && (row * 640 + col) <= 64639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 64640 && (row * 640 + col) <= 64679) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 64680 && (row * 640 + col) <= 65038) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 65039 && (row * 640 + col) <= 65041) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65042 && (row * 640 + col) <= 65089) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 65090 && (row * 640 + col) <= 65118) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65119 && (row * 640 + col) <= 65678) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 65679 && (row * 640 + col) <= 65681) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 65682 && (row * 640 + col) <= 65725) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 65726 && (row * 640 + col) <= 65763) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 65764 && (row * 640 + col) <= 66318) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 66319 && (row * 640 + col) <= 66321) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66322 && (row * 640 + col) <= 66364) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 66365 && (row * 640 + col) <= 66404) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 66405 && (row * 640 + col) <= 66958) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 66959 && (row * 640 + col) <= 66961) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 66962 && (row * 640 + col) <= 67004) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 67005 && (row * 640 + col) <= 67044) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67045 && (row * 640 + col) <= 67593) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 67594 && (row * 640 + col) <= 67606) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 67607 && (row * 640 + col) <= 67642) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 67643 && (row * 640 + col) <= 67686) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 67687 && (row * 640 + col) <= 68232) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 68233 && (row * 640 + col) <= 68246) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68247 && (row * 640 + col) <= 68281) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 68282 && (row * 640 + col) <= 68327) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68328 && (row * 640 + col) <= 68872) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 68873 && (row * 640 + col) <= 68887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 68888 && (row * 640 + col) <= 68921) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 68922 && (row * 640 + col) <= 68967) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 68968 && (row * 640 + col) <= 69512) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 69513 && (row * 640 + col) <= 69527) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 69528 && (row * 640 + col) <= 69558) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 69559 && (row * 640 + col) <= 69607) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 69608 && (row * 640 + col) <= 70152) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 70153 && (row * 640 + col) <= 70166) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70167 && (row * 640 + col) <= 70198) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 70199 && (row * 640 + col) <= 70247) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70248 && (row * 640 + col) <= 70792) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 70793 && (row * 640 + col) <= 70807) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 70808 && (row * 640 + col) <= 70838) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 70839 && (row * 640 + col) <= 70887) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 70888 && (row * 640 + col) <= 71426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 71427 && (row * 640 + col) <= 71452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 71453 && (row * 640 + col) <= 71476) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 71477 && (row * 640 + col) <= 71529) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 71530 && (row * 640 + col) <= 72066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 72067 && (row * 640 + col) <= 72092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72093 && (row * 640 + col) <= 72115) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 72116 && (row * 640 + col) <= 72170) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72171 && (row * 640 + col) <= 72706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 72707 && (row * 640 + col) <= 72732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 72733 && (row * 640 + col) <= 72755) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 72756 && (row * 640 + col) <= 72810) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 72811 && (row * 640 + col) <= 73346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 73347 && (row * 640 + col) <= 73372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 73373 && (row * 640 + col) <= 73387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 73388 && (row * 640 + col) <= 73450) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 73451 && (row * 640 + col) <= 73986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 73987 && (row * 640 + col) <= 74012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74013 && (row * 640 + col) <= 74026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 74027 && (row * 640 + col) <= 74090) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74091 && (row * 640 + col) <= 74626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 74627 && (row * 640 + col) <= 74652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 74653 && (row * 640 + col) <= 74666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 74667 && (row * 640 + col) <= 74730) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 74731 && (row * 640 + col) <= 75266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 75267 && (row * 640 + col) <= 75292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75293 && (row * 640 + col) <= 75301) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 75302 && (row * 640 + col) <= 75370) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 75371 && (row * 640 + col) <= 75906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 75907 && (row * 640 + col) <= 75932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 75933 && (row * 640 + col) <= 75941) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 75942 && (row * 640 + col) <= 76010) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76011 && (row * 640 + col) <= 76546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 76547 && (row * 640 + col) <= 76572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 76573 && (row * 640 + col) <= 76580) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 76581 && (row * 640 + col) <= 76650) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 76651 && (row * 640 + col) <= 77186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 77187 && (row * 640 + col) <= 77212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77213 && (row * 640 + col) <= 77218) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 77219 && (row * 640 + col) <= 77295) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77296 && (row * 640 + col) <= 77826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 77827 && (row * 640 + col) <= 77852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 77853 && (row * 640 + col) <= 77858) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 77859 && (row * 640 + col) <= 77936) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 77937 && (row * 640 + col) <= 78466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 78467 && (row * 640 + col) <= 78492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 78493 && (row * 640 + col) <= 78498) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 78499 && (row * 640 + col) <= 78577) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 78578 && (row * 640 + col) <= 79106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 79107 && (row * 640 + col) <= 79132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79133 && (row * 640 + col) <= 79138) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 79139 && (row * 640 + col) <= 79218) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79219 && (row * 640 + col) <= 79746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 79747 && (row * 640 + col) <= 79772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 79773 && (row * 640 + col) <= 79778) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 79779 && (row * 640 + col) <= 79858) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 79859 && (row * 640 + col) <= 80386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 80387 && (row * 640 + col) <= 80412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 80413 && (row * 640 + col) <= 80416) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 80417 && (row * 640 + col) <= 80503) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 80504 && (row * 640 + col) <= 81026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 81027 && (row * 640 + col) <= 81052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81053 && (row * 640 + col) <= 81055) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 81056 && (row * 640 + col) <= 81144) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81145 && (row * 640 + col) <= 81666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 81667 && (row * 640 + col) <= 81692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 81693 && (row * 640 + col) <= 81695) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 81696 && (row * 640 + col) <= 81784) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 81785 && (row * 640 + col) <= 82306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 82307 && (row * 640 + col) <= 82332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82333 && (row * 640 + col) <= 82333) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 82334 && (row * 640 + col) <= 82426) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 82427 && (row * 640 + col) <= 82946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 82947 && (row * 640 + col) <= 82972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 82973 && (row * 640 + col) <= 83067) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83068 && (row * 640 + col) <= 83586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 83587 && (row * 640 + col) <= 83612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 83613 && (row * 640 + col) <= 83707) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 83708 && (row * 640 + col) <= 84226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 84227 && (row * 640 + col) <= 84252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84253 && (row * 640 + col) <= 84352) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84353 && (row * 640 + col) <= 84866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 84867 && (row * 640 + col) <= 84892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 84893 && (row * 640 + col) <= 84993) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 84994 && (row * 640 + col) <= 85506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 85507 && (row * 640 + col) <= 85532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 85533 && (row * 640 + col) <= 85632) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 85633 && (row * 640 + col) <= 86146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 86147 && (row * 640 + col) <= 86172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86173 && (row * 640 + col) <= 86190) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86191 && (row * 640 + col) <= 86204) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 86205 && (row * 640 + col) <= 86258) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86259 && (row * 640 + col) <= 86786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 86787 && (row * 640 + col) <= 86812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 86813 && (row * 640 + col) <= 86829) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86830 && (row * 640 + col) <= 86844) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 86845 && (row * 640 + col) <= 86898) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 86899 && (row * 640 + col) <= 87426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87427 && (row * 640 + col) <= 87452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 87453 && (row * 640 + col) <= 87453) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87454 && (row * 640 + col) <= 87469) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87470 && (row * 640 + col) <= 87484) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87485 && (row * 640 + col) <= 87488) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87489 && (row * 640 + col) <= 87490) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87491 && (row * 640 + col) <= 87502) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87503 && (row * 640 + col) <= 87504) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87505 && (row * 640 + col) <= 87513) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87514 && (row * 640 + col) <= 87517) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 87518 && (row * 640 + col) <= 87538) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 87539 && (row * 640 + col) <= 88066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88067 && (row * 640 + col) <= 88092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88093 && (row * 640 + col) <= 88101) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88102 && (row * 640 + col) <= 88103) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88104 && (row * 640 + col) <= 88125) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88126 && (row * 640 + col) <= 88126) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88127 && (row * 640 + col) <= 88136) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88137 && (row * 640 + col) <= 88138) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88139 && (row * 640 + col) <= 88147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88148 && (row * 640 + col) <= 88149) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88150 && (row * 640 + col) <= 88159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88160 && (row * 640 + col) <= 88160) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88161 && (row * 640 + col) <= 88170) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88171 && (row * 640 + col) <= 88172) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 88173 && (row * 640 + col) <= 88706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 88707 && (row * 640 + col) <= 88732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 88733 && (row * 640 + col) <= 89346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 89347 && (row * 640 + col) <= 89372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89373 && (row * 640 + col) <= 89946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 89947 && (row * 640 + col) <= 89966) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 89967 && (row * 640 + col) <= 89986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 89987 && (row * 640 + col) <= 90012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90013 && (row * 640 + col) <= 90586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 90587 && (row * 640 + col) <= 90606) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90607 && (row * 640 + col) <= 90626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 90627 && (row * 640 + col) <= 90652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 90653 && (row * 640 + col) <= 91226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 91227 && (row * 640 + col) <= 91246) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91247 && (row * 640 + col) <= 91266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 91267 && (row * 640 + col) <= 91292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91293 && (row * 640 + col) <= 91866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 91867 && (row * 640 + col) <= 91886) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91887 && (row * 640 + col) <= 91906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 91907 && (row * 640 + col) <= 91932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 91933 && (row * 640 + col) <= 92506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 92507 && (row * 640 + col) <= 92526) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 92527 && (row * 640 + col) <= 92546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 92547 && (row * 640 + col) <= 92572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 92573 && (row * 640 + col) <= 93146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 93147 && (row * 640 + col) <= 93166) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 93167 && (row * 640 + col) <= 93186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 93187 && (row * 640 + col) <= 93212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 93213 && (row * 640 + col) <= 93437) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 93438 && (row * 640 + col) <= 93439) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 93440 && (row * 640 + col) <= 93786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 93787 && (row * 640 + col) <= 93806) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 93807 && (row * 640 + col) <= 93826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 93827 && (row * 640 + col) <= 93852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 93853 && (row * 640 + col) <= 94076) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 94077 && (row * 640 + col) <= 94079) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94080 && (row * 640 + col) <= 94426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 94427 && (row * 640 + col) <= 94446) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 94447 && (row * 640 + col) <= 94466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 94467 && (row * 640 + col) <= 94492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 94493 && (row * 640 + col) <= 94716) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 94717 && (row * 640 + col) <= 94719) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 94720 && (row * 640 + col) <= 95066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 95067 && (row * 640 + col) <= 95086) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 95087 && (row * 640 + col) <= 95107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 95108 && (row * 640 + col) <= 95132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 95133 && (row * 640 + col) <= 95354) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 95355 && (row * 640 + col) <= 95359) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 95360 && (row * 640 + col) <= 95706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 95707 && (row * 640 + col) <= 95726) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 95727 && (row * 640 + col) <= 95747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 95748 && (row * 640 + col) <= 95772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 95773 && (row * 640 + col) <= 95992) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 95993 && (row * 640 + col) <= 95999) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96000 && (row * 640 + col) <= 96103) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96104 && (row * 640 + col) <= 96105) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96106 && (row * 640 + col) <= 96109) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96110 && (row * 640 + col) <= 96110) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96111 && (row * 640 + col) <= 96120) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96121 && (row * 640 + col) <= 96122) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96123 && (row * 640 + col) <= 96126) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96127 && (row * 640 + col) <= 96127) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96128 && (row * 640 + col) <= 96131) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96132 && (row * 640 + col) <= 96133) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96134 && (row * 640 + col) <= 96137) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96138 && (row * 640 + col) <= 96139) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96140 && (row * 640 + col) <= 96346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96347 && (row * 640 + col) <= 96366) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 96367 && (row * 640 + col) <= 96387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96388 && (row * 640 + col) <= 96412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 96413 && (row * 640 + col) <= 96631) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96632 && (row * 640 + col) <= 96639) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96640 && (row * 640 + col) <= 96676) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 96677 && (row * 640 + col) <= 96742) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96743 && (row * 640 + col) <= 96753) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96754 && (row * 640 + col) <= 96759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96760 && (row * 640 + col) <= 96780) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 96781 && (row * 640 + col) <= 96880) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96881 && (row * 640 + col) <= 96883) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 96884 && (row * 640 + col) <= 96946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96947 && (row * 640 + col) <= 96974) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 96975 && (row * 640 + col) <= 96986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 96987 && (row * 640 + col) <= 97006) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97007 && (row * 640 + col) <= 97026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97027 && (row * 640 + col) <= 97052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97053 && (row * 640 + col) <= 97144) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97145 && (row * 640 + col) <= 97167) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97168 && (row * 640 + col) <= 97268) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97269 && (row * 640 + col) <= 97279) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97280 && (row * 640 + col) <= 97316) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97317 && (row * 640 + col) <= 97381) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97382 && (row * 640 + col) <= 97394) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97395 && (row * 640 + col) <= 97398) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97399 && (row * 640 + col) <= 97420) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97421 && (row * 640 + col) <= 97520) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97521 && (row * 640 + col) <= 97523) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97524 && (row * 640 + col) <= 97586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97587 && (row * 640 + col) <= 97615) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97616 && (row * 640 + col) <= 97626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97627 && (row * 640 + col) <= 97646) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97647 && (row * 640 + col) <= 97666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97667 && (row * 640 + col) <= 97692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97693 && (row * 640 + col) <= 97784) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97785 && (row * 640 + col) <= 97807) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97808 && (row * 640 + col) <= 97907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 97908 && (row * 640 + col) <= 97919) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 97920 && (row * 640 + col) <= 97956) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 97957 && (row * 640 + col) <= 98020) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98021 && (row * 640 + col) <= 98034) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98035 && (row * 640 + col) <= 98038) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98039 && (row * 640 + col) <= 98061) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98062 && (row * 640 + col) <= 98160) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98161 && (row * 640 + col) <= 98163) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98164 && (row * 640 + col) <= 98226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98227 && (row * 640 + col) <= 98255) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98256 && (row * 640 + col) <= 98266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98267 && (row * 640 + col) <= 98286) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98287 && (row * 640 + col) <= 98306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98307 && (row * 640 + col) <= 98332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98333 && (row * 640 + col) <= 98424) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98425 && (row * 640 + col) <= 98447) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98448 && (row * 640 + col) <= 98547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98548 && (row * 640 + col) <= 98559) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98560 && (row * 640 + col) <= 98596) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98597 && (row * 640 + col) <= 98656) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98657 && (row * 640 + col) <= 98703) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 98704 && (row * 640 + col) <= 98731) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98732 && (row * 640 + col) <= 98757) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98758 && (row * 640 + col) <= 98780) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98781 && (row * 640 + col) <= 98783) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98784 && (row * 640 + col) <= 98800) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98801 && (row * 640 + col) <= 98803) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98804 && (row * 640 + col) <= 98866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98867 && (row * 640 + col) <= 98895) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98896 && (row * 640 + col) <= 98906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98907 && (row * 640 + col) <= 98926) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98927 && (row * 640 + col) <= 98947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 98948 && (row * 640 + col) <= 98972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 98973 && (row * 640 + col) <= 99064) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99065 && (row * 640 + col) <= 99087) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99088 && (row * 640 + col) <= 99181) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99182 && (row * 640 + col) <= 99199) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99200 && (row * 640 + col) <= 99236) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99237 && (row * 640 + col) <= 99296) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99297 && (row * 640 + col) <= 99343) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99344 && (row * 640 + col) <= 99371) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99372 && (row * 640 + col) <= 99397) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99398 && (row * 640 + col) <= 99420) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99421 && (row * 640 + col) <= 99423) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99424 && (row * 640 + col) <= 99440) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99441 && (row * 640 + col) <= 99443) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99444 && (row * 640 + col) <= 99506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99507 && (row * 640 + col) <= 99535) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99536 && (row * 640 + col) <= 99546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99547 && (row * 640 + col) <= 99566) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99567 && (row * 640 + col) <= 99587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99588 && (row * 640 + col) <= 99612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99613 && (row * 640 + col) <= 99704) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99705 && (row * 640 + col) <= 99727) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99728 && (row * 640 + col) <= 99820) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99821 && (row * 640 + col) <= 99839) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99840 && (row * 640 + col) <= 99876) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 99877 && (row * 640 + col) <= 99934) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 99935 && (row * 640 + col) <= 99984) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 99985 && (row * 640 + col) <= 100011) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100012 && (row * 640 + col) <= 100037) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100038 && (row * 640 + col) <= 100060) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100061 && (row * 640 + col) <= 100063) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100064 && (row * 640 + col) <= 100080) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100081 && (row * 640 + col) <= 100083) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100084 && (row * 640 + col) <= 100146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100147 && (row * 640 + col) <= 100175) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100176 && (row * 640 + col) <= 100186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100187 && (row * 640 + col) <= 100206) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100207 && (row * 640 + col) <= 100227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100228 && (row * 640 + col) <= 100252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100253 && (row * 640 + col) <= 100344) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100345 && (row * 640 + col) <= 100367) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100368 && (row * 640 + col) <= 100450) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100451 && (row * 640 + col) <= 100456) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100457 && (row * 640 + col) <= 100459) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100460 && (row * 640 + col) <= 100479) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100480 && (row * 640 + col) <= 100516) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100517 && (row * 640 + col) <= 100573) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100574 && (row * 640 + col) <= 100623) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 100624 && (row * 640 + col) <= 100651) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100652 && (row * 640 + col) <= 100677) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100678 && (row * 640 + col) <= 100700) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100701 && (row * 640 + col) <= 100703) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100704 && (row * 640 + col) <= 100717) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100718 && (row * 640 + col) <= 100725) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100726 && (row * 640 + col) <= 100786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100787 && (row * 640 + col) <= 100815) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100816 && (row * 640 + col) <= 100826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100827 && (row * 640 + col) <= 100852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100853 && (row * 640 + col) <= 100867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100868 && (row * 640 + col) <= 100892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100893 && (row * 640 + col) <= 100961) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100962 && (row * 640 + col) <= 100978) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 100979 && (row * 640 + col) <= 100984) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 100985 && (row * 640 + col) <= 101007) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101008 && (row * 640 + col) <= 101089) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101090 && (row * 640 + col) <= 101119) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101120 && (row * 640 + col) <= 101156) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101157 && (row * 640 + col) <= 101212) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101213 && (row * 640 + col) <= 101263) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101264 && (row * 640 + col) <= 101291) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101292 && (row * 640 + col) <= 101317) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101318 && (row * 640 + col) <= 101340) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101341 && (row * 640 + col) <= 101343) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101344 && (row * 640 + col) <= 101357) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101358 && (row * 640 + col) <= 101366) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101367 && (row * 640 + col) <= 101426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101427 && (row * 640 + col) <= 101455) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101456 && (row * 640 + col) <= 101466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101467 && (row * 640 + col) <= 101492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101493 && (row * 640 + col) <= 101507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101508 && (row * 640 + col) <= 101532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101533 && (row * 640 + col) <= 101601) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101602 && (row * 640 + col) <= 101618) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101619 && (row * 640 + col) <= 101624) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101625 && (row * 640 + col) <= 101647) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101648 && (row * 640 + col) <= 101729) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101730 && (row * 640 + col) <= 101759) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101760 && (row * 640 + col) <= 101796) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101797 && (row * 640 + col) <= 101850) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101851 && (row * 640 + col) <= 101904) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 101905 && (row * 640 + col) <= 101931) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101932 && (row * 640 + col) <= 101957) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101958 && (row * 640 + col) <= 101980) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101981 && (row * 640 + col) <= 101983) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 101984 && (row * 640 + col) <= 101997) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 101998 && (row * 640 + col) <= 102006) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102007 && (row * 640 + col) <= 102066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102067 && (row * 640 + col) <= 102095) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102096 && (row * 640 + col) <= 102106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102107 && (row * 640 + col) <= 102132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102133 && (row * 640 + col) <= 102147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102148 && (row * 640 + col) <= 102172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102173 && (row * 640 + col) <= 102241) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102242 && (row * 640 + col) <= 102258) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102259 && (row * 640 + col) <= 102264) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102265 && (row * 640 + col) <= 102287) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102288 && (row * 640 + col) <= 102362) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102363 && (row * 640 + col) <= 102399) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102400 && (row * 640 + col) <= 102436) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102437 && (row * 640 + col) <= 102490) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102491 && (row * 640 + col) <= 102543) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 102544 && (row * 640 + col) <= 102571) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102572 && (row * 640 + col) <= 102597) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102598 && (row * 640 + col) <= 102620) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102621 && (row * 640 + col) <= 102623) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102624 && (row * 640 + col) <= 102637) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102638 && (row * 640 + col) <= 102646) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102647 && (row * 640 + col) <= 102669) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102670 && (row * 640 + col) <= 102691) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102692 && (row * 640 + col) <= 102706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102707 && (row * 640 + col) <= 102735) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102736 && (row * 640 + col) <= 102746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102747 && (row * 640 + col) <= 102772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102773 && (row * 640 + col) <= 102787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102788 && (row * 640 + col) <= 102812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102813 && (row * 640 + col) <= 102881) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102882 && (row * 640 + col) <= 102898) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102899 && (row * 640 + col) <= 102904) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 102905 && (row * 640 + col) <= 102927) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 102928 && (row * 640 + col) <= 103001) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103002 && (row * 640 + col) <= 103039) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103040 && (row * 640 + col) <= 103076) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103077 && (row * 640 + col) <= 103129) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103130 && (row * 640 + col) <= 103183) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103184 && (row * 640 + col) <= 103211) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103212 && (row * 640 + col) <= 103237) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103238 && (row * 640 + col) <= 103260) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103261 && (row * 640 + col) <= 103263) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103264 && (row * 640 + col) <= 103277) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103278 && (row * 640 + col) <= 103286) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103287 && (row * 640 + col) <= 103309) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103310 && (row * 640 + col) <= 103331) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103332 && (row * 640 + col) <= 103346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103347 && (row * 640 + col) <= 103375) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103376 && (row * 640 + col) <= 103386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103387 && (row * 640 + col) <= 103412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103413 && (row * 640 + col) <= 103427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103428 && (row * 640 + col) <= 103452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103453 && (row * 640 + col) <= 103521) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103522 && (row * 640 + col) <= 103538) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103539 && (row * 640 + col) <= 103544) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103545 && (row * 640 + col) <= 103567) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103568 && (row * 640 + col) <= 103638) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103639 && (row * 640 + col) <= 103639) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103640 && (row * 640 + col) <= 103640) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103641 && (row * 640 + col) <= 103679) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103680 && (row * 640 + col) <= 103716) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103717 && (row * 640 + col) <= 103767) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103768 && (row * 640 + col) <= 103823) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 103824 && (row * 640 + col) <= 103851) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103852 && (row * 640 + col) <= 103877) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103878 && (row * 640 + col) <= 103900) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103901 && (row * 640 + col) <= 103903) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103904 && (row * 640 + col) <= 103917) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103918 && (row * 640 + col) <= 103926) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103927 && (row * 640 + col) <= 103949) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103950 && (row * 640 + col) <= 103971) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 103972 && (row * 640 + col) <= 103986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 103987 && (row * 640 + col) <= 104015) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104016 && (row * 640 + col) <= 104026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104027 && (row * 640 + col) <= 104052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104053 && (row * 640 + col) <= 104067) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104068 && (row * 640 + col) <= 104092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104093 && (row * 640 + col) <= 104161) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104162 && (row * 640 + col) <= 104178) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104179 && (row * 640 + col) <= 104184) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104185 && (row * 640 + col) <= 104207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104208 && (row * 640 + col) <= 104273) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104274 && (row * 640 + col) <= 104319) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104320 && (row * 640 + col) <= 104356) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104357 && (row * 640 + col) <= 104407) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104408 && (row * 640 + col) <= 104463) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104464 && (row * 640 + col) <= 104491) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104492 && (row * 640 + col) <= 104517) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104518 && (row * 640 + col) <= 104540) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104541 && (row * 640 + col) <= 104543) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104544 && (row * 640 + col) <= 104555) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104556 && (row * 640 + col) <= 104568) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104569 && (row * 640 + col) <= 104589) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104590 && (row * 640 + col) <= 104611) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104612 && (row * 640 + col) <= 104626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104627 && (row * 640 + col) <= 104655) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104656 && (row * 640 + col) <= 104666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104667 && (row * 640 + col) <= 104692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104693 && (row * 640 + col) <= 104707) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104708 && (row * 640 + col) <= 104732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104733 && (row * 640 + col) <= 104801) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104802 && (row * 640 + col) <= 104818) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104819 && (row * 640 + col) <= 104824) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104825 && (row * 640 + col) <= 104847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104848 && (row * 640 + col) <= 104912) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 104913 && (row * 640 + col) <= 104959) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 104960 && (row * 640 + col) <= 104996) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 104997 && (row * 640 + col) <= 105047) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105048 && (row * 640 + col) <= 105104) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105105 && (row * 640 + col) <= 105131) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105132 && (row * 640 + col) <= 105157) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105158 && (row * 640 + col) <= 105180) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105181 && (row * 640 + col) <= 105183) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105184 && (row * 640 + col) <= 105195) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105196 && (row * 640 + col) <= 105208) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105209 && (row * 640 + col) <= 105229) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105230 && (row * 640 + col) <= 105251) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105252 && (row * 640 + col) <= 105266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105267 && (row * 640 + col) <= 105295) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105296 && (row * 640 + col) <= 105306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105307 && (row * 640 + col) <= 105332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105333 && (row * 640 + col) <= 105347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105348 && (row * 640 + col) <= 105372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105373 && (row * 640 + col) <= 105441) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105442 && (row * 640 + col) <= 105458) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105459 && (row * 640 + col) <= 105464) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105465 && (row * 640 + col) <= 105487) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105488 && (row * 640 + col) <= 105552) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105553 && (row * 640 + col) <= 105599) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105600 && (row * 640 + col) <= 105636) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105637 && (row * 640 + col) <= 105687) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105688 && (row * 640 + col) <= 105745) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 105746 && (row * 640 + col) <= 105771) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105772 && (row * 640 + col) <= 105797) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105798 && (row * 640 + col) <= 105820) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105821 && (row * 640 + col) <= 105823) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105824 && (row * 640 + col) <= 105835) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105836 && (row * 640 + col) <= 105848) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105849 && (row * 640 + col) <= 105869) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105870 && (row * 640 + col) <= 105891) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105892 && (row * 640 + col) <= 105906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105907 && (row * 640 + col) <= 105935) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105936 && (row * 640 + col) <= 105946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105947 && (row * 640 + col) <= 105972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 105973 && (row * 640 + col) <= 105987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 105988 && (row * 640 + col) <= 106012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106013 && (row * 640 + col) <= 106081) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106082 && (row * 640 + col) <= 106098) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106099 && (row * 640 + col) <= 106104) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106105 && (row * 640 + col) <= 106127) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106128 && (row * 640 + col) <= 106190) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106191 && (row * 640 + col) <= 106239) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106240 && (row * 640 + col) <= 106276) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106277 && (row * 640 + col) <= 106327) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106328 && (row * 640 + col) <= 106386) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106387 && (row * 640 + col) <= 106411) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106412 && (row * 640 + col) <= 106437) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106438 && (row * 640 + col) <= 106457) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106458 && (row * 640 + col) <= 106465) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106466 && (row * 640 + col) <= 106475) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106476 && (row * 640 + col) <= 106488) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106489 && (row * 640 + col) <= 106509) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106510 && (row * 640 + col) <= 106531) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106532 && (row * 640 + col) <= 106546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106547 && (row * 640 + col) <= 106575) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106576 && (row * 640 + col) <= 106586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106587 && (row * 640 + col) <= 106612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106613 && (row * 640 + col) <= 106627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106628 && (row * 640 + col) <= 106652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106653 && (row * 640 + col) <= 106721) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106722 && (row * 640 + col) <= 106738) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106739 && (row * 640 + col) <= 106744) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106745 && (row * 640 + col) <= 106767) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106768 && (row * 640 + col) <= 106829) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106830 && (row * 640 + col) <= 106879) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 106880 && (row * 640 + col) <= 106916) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 106917 && (row * 640 + col) <= 106966) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 106967 && (row * 640 + col) <= 107027) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107028 && (row * 640 + col) <= 107051) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107052 && (row * 640 + col) <= 107077) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107078 && (row * 640 + col) <= 107097) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107098 && (row * 640 + col) <= 107105) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107106 && (row * 640 + col) <= 107115) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107116 && (row * 640 + col) <= 107128) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107129 && (row * 640 + col) <= 107149) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107150 && (row * 640 + col) <= 107171) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107172 && (row * 640 + col) <= 107186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107187 && (row * 640 + col) <= 107215) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107216 && (row * 640 + col) <= 107226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107227 && (row * 640 + col) <= 107252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107253 && (row * 640 + col) <= 107267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107268 && (row * 640 + col) <= 107292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107293 && (row * 640 + col) <= 107361) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107362 && (row * 640 + col) <= 107378) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107379 && (row * 640 + col) <= 107384) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107385 && (row * 640 + col) <= 107407) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107408 && (row * 640 + col) <= 107469) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107470 && (row * 640 + col) <= 107519) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107520 && (row * 640 + col) <= 107556) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107557 && (row * 640 + col) <= 107605) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107606 && (row * 640 + col) <= 107669) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 107670 && (row * 640 + col) <= 107691) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107692 && (row * 640 + col) <= 107717) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107718 && (row * 640 + col) <= 107737) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107738 && (row * 640 + col) <= 107745) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107746 && (row * 640 + col) <= 107755) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107756 && (row * 640 + col) <= 107768) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107769 && (row * 640 + col) <= 107789) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107790 && (row * 640 + col) <= 107811) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107812 && (row * 640 + col) <= 107826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107827 && (row * 640 + col) <= 107855) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107856 && (row * 640 + col) <= 107866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107867 && (row * 640 + col) <= 107892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107893 && (row * 640 + col) <= 107907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 107908 && (row * 640 + col) <= 107932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 107933 && (row * 640 + col) <= 108001) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108002 && (row * 640 + col) <= 108018) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108019 && (row * 640 + col) <= 108024) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108025 && (row * 640 + col) <= 108047) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108048 && (row * 640 + col) <= 108104) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108105 && (row * 640 + col) <= 108159) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108160 && (row * 640 + col) <= 108196) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108197 && (row * 640 + col) <= 108244) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108245 && (row * 640 + col) <= 108309) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108310 && (row * 640 + col) <= 108331) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108332 && (row * 640 + col) <= 108357) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108358 && (row * 640 + col) <= 108363) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108364 && (row * 640 + col) <= 108385) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108386 && (row * 640 + col) <= 108395) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108396 && (row * 640 + col) <= 108408) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108409 && (row * 640 + col) <= 108429) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108430 && (row * 640 + col) <= 108451) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108452 && (row * 640 + col) <= 108466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108467 && (row * 640 + col) <= 108495) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108496 && (row * 640 + col) <= 108506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108507 && (row * 640 + col) <= 108532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108533 && (row * 640 + col) <= 108547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108548 && (row * 640 + col) <= 108572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108573 && (row * 640 + col) <= 108641) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108642 && (row * 640 + col) <= 108658) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108659 && (row * 640 + col) <= 108664) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108665 && (row * 640 + col) <= 108687) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108688 && (row * 640 + col) <= 108743) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108744 && (row * 640 + col) <= 108777) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108778 && (row * 640 + col) <= 108786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108787 && (row * 640 + col) <= 108799) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108800 && (row * 640 + col) <= 108836) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108837 && (row * 640 + col) <= 108882) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108883 && (row * 640 + col) <= 108949) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108950 && (row * 640 + col) <= 108952) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108953 && (row * 640 + col) <= 108954) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 108955 && (row * 640 + col) <= 108971) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 108972 && (row * 640 + col) <= 108997) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 108998 && (row * 640 + col) <= 109003) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109004 && (row * 640 + col) <= 109025) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109026 && (row * 640 + col) <= 109035) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109036 && (row * 640 + col) <= 109048) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109049 && (row * 640 + col) <= 109069) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109070 && (row * 640 + col) <= 109091) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109092 && (row * 640 + col) <= 109106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109107 && (row * 640 + col) <= 109135) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109136 && (row * 640 + col) <= 109146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109147 && (row * 640 + col) <= 109172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109173 && (row * 640 + col) <= 109187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109188 && (row * 640 + col) <= 109212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109213 && (row * 640 + col) <= 109281) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109282 && (row * 640 + col) <= 109298) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109299 && (row * 640 + col) <= 109304) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109305 && (row * 640 + col) <= 109327) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109328 && (row * 640 + col) <= 109383) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109384 && (row * 640 + col) <= 109417) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109418 && (row * 640 + col) <= 109427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109428 && (row * 640 + col) <= 109439) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109440 && (row * 640 + col) <= 109477) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109478 && (row * 640 + col) <= 109522) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109523 && (row * 640 + col) <= 109595) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 109596 && (row * 640 + col) <= 109611) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109612 && (row * 640 + col) <= 109637) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109638 && (row * 640 + col) <= 109643) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109644 && (row * 640 + col) <= 109666) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109667 && (row * 640 + col) <= 109675) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109676 && (row * 640 + col) <= 109688) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109689 && (row * 640 + col) <= 109709) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109710 && (row * 640 + col) <= 109731) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109732 && (row * 640 + col) <= 109746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109747 && (row * 640 + col) <= 109775) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109776 && (row * 640 + col) <= 109786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109787 && (row * 640 + col) <= 109812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109813 && (row * 640 + col) <= 109827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109828 && (row * 640 + col) <= 109852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109853 && (row * 640 + col) <= 109921) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109922 && (row * 640 + col) <= 109938) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109939 && (row * 640 + col) <= 109944) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 109945 && (row * 640 + col) <= 109967) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 109968 && (row * 640 + col) <= 110024) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110025 && (row * 640 + col) <= 110056) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110057 && (row * 640 + col) <= 110067) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110068 && (row * 640 + col) <= 110079) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110080 && (row * 640 + col) <= 110125) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110126 && (row * 640 + col) <= 110161) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110162 && (row * 640 + col) <= 110217) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110218 && (row * 640 + col) <= 110231) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110232 && (row * 640 + col) <= 110235) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110236 && (row * 640 + col) <= 110251) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110252 && (row * 640 + col) <= 110277) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110278 && (row * 640 + col) <= 110283) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110284 && (row * 640 + col) <= 110308) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110309 && (row * 640 + col) <= 110315) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110316 && (row * 640 + col) <= 110328) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110329 && (row * 640 + col) <= 110349) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110350 && (row * 640 + col) <= 110371) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110372 && (row * 640 + col) <= 110386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110387 && (row * 640 + col) <= 110415) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110416 && (row * 640 + col) <= 110426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110427 && (row * 640 + col) <= 110452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110453 && (row * 640 + col) <= 110467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110468 && (row * 640 + col) <= 110492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110493 && (row * 640 + col) <= 110561) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110562 && (row * 640 + col) <= 110578) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110579 && (row * 640 + col) <= 110584) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110585 && (row * 640 + col) <= 110607) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110608 && (row * 640 + col) <= 110664) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110665 && (row * 640 + col) <= 110666) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110667 && (row * 640 + col) <= 110709) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110710 && (row * 640 + col) <= 110710) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110711 && (row * 640 + col) <= 110719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110720 && (row * 640 + col) <= 110765) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110766 && (row * 640 + col) <= 110796) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110797 && (row * 640 + col) <= 110857) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110858 && (row * 640 + col) <= 110871) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110872 && (row * 640 + col) <= 110875) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 110876 && (row * 640 + col) <= 110891) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110892 && (row * 640 + col) <= 110917) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110918 && (row * 640 + col) <= 110923) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110924 && (row * 640 + col) <= 110948) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110949 && (row * 640 + col) <= 110955) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110956 && (row * 640 + col) <= 110968) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 110969 && (row * 640 + col) <= 110989) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 110990 && (row * 640 + col) <= 111011) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111012 && (row * 640 + col) <= 111026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111027 && (row * 640 + col) <= 111055) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111056 && (row * 640 + col) <= 111066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111067 && (row * 640 + col) <= 111092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111093 && (row * 640 + col) <= 111107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111108 && (row * 640 + col) <= 111132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111133 && (row * 640 + col) <= 111201) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111202 && (row * 640 + col) <= 111218) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111219 && (row * 640 + col) <= 111224) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111225 && (row * 640 + col) <= 111247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111248 && (row * 640 + col) <= 111359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111360 && (row * 640 + col) <= 111405) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111406 && (row * 640 + col) <= 111435) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111436 && (row * 640 + col) <= 111497) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 111498 && (row * 640 + col) <= 111588) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111589 && (row * 640 + col) <= 111595) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111596 && (row * 640 + col) <= 111608) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111609 && (row * 640 + col) <= 111629) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111630 && (row * 640 + col) <= 111651) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111652 && (row * 640 + col) <= 111666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111667 && (row * 640 + col) <= 111695) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111696 && (row * 640 + col) <= 111706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111707 && (row * 640 + col) <= 111732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111733 && (row * 640 + col) <= 111747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111748 && (row * 640 + col) <= 111772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111773 && (row * 640 + col) <= 111841) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111842 && (row * 640 + col) <= 111858) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111859 && (row * 640 + col) <= 111864) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 111865 && (row * 640 + col) <= 111887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 111888 && (row * 640 + col) <= 111999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112000 && (row * 640 + col) <= 112045) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112046 && (row * 640 + col) <= 112075) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112076 && (row * 640 + col) <= 112137) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112138 && (row * 640 + col) <= 112228) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112229 && (row * 640 + col) <= 112235) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112236 && (row * 640 + col) <= 112248) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112249 && (row * 640 + col) <= 112269) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112270 && (row * 640 + col) <= 112291) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112292 && (row * 640 + col) <= 112306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112307 && (row * 640 + col) <= 112335) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112336 && (row * 640 + col) <= 112346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112347 && (row * 640 + col) <= 112372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112373 && (row * 640 + col) <= 112387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112388 && (row * 640 + col) <= 112412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112413 && (row * 640 + col) <= 112481) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112482 && (row * 640 + col) <= 112498) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112499 && (row * 640 + col) <= 112504) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112505 && (row * 640 + col) <= 112527) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112528 && (row * 640 + col) <= 112639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112640 && (row * 640 + col) <= 112685) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112686 && (row * 640 + col) <= 112714) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112715 && (row * 640 + col) <= 112777) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 112778 && (row * 640 + col) <= 112868) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112869 && (row * 640 + col) <= 112875) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112876 && (row * 640 + col) <= 112888) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112889 && (row * 640 + col) <= 112909) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112910 && (row * 640 + col) <= 112931) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112932 && (row * 640 + col) <= 112946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112947 && (row * 640 + col) <= 112975) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 112976 && (row * 640 + col) <= 112986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 112987 && (row * 640 + col) <= 113012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113013 && (row * 640 + col) <= 113027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113028 && (row * 640 + col) <= 113052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113053 && (row * 640 + col) <= 113121) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113122 && (row * 640 + col) <= 113138) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113139 && (row * 640 + col) <= 113144) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113145 && (row * 640 + col) <= 113167) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113168 && (row * 640 + col) <= 113279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113280 && (row * 640 + col) <= 113325) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113326 && (row * 640 + col) <= 113350) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113351 && (row * 640 + col) <= 113417) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 113418 && (row * 640 + col) <= 113508) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113509 && (row * 640 + col) <= 113515) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113516 && (row * 640 + col) <= 113528) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113529 && (row * 640 + col) <= 113549) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113550 && (row * 640 + col) <= 113571) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113572 && (row * 640 + col) <= 113586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113587 && (row * 640 + col) <= 113615) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113616 && (row * 640 + col) <= 113626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113627 && (row * 640 + col) <= 113652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113653 && (row * 640 + col) <= 113667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113668 && (row * 640 + col) <= 113692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113693 && (row * 640 + col) <= 113761) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113762 && (row * 640 + col) <= 113778) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113779 && (row * 640 + col) <= 113784) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113785 && (row * 640 + col) <= 113807) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113808 && (row * 640 + col) <= 113919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113920 && (row * 640 + col) <= 113965) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 113966 && (row * 640 + col) <= 113990) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 113991 && (row * 640 + col) <= 114057) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114058 && (row * 640 + col) <= 114148) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114149 && (row * 640 + col) <= 114155) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114156 && (row * 640 + col) <= 114168) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114169 && (row * 640 + col) <= 114189) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114190 && (row * 640 + col) <= 114211) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114212 && (row * 640 + col) <= 114226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114227 && (row * 640 + col) <= 114255) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114256 && (row * 640 + col) <= 114266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114267 && (row * 640 + col) <= 114292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114293 && (row * 640 + col) <= 114307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114308 && (row * 640 + col) <= 114332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114333 && (row * 640 + col) <= 114401) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114402 && (row * 640 + col) <= 114418) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114419 && (row * 640 + col) <= 114424) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114425 && (row * 640 + col) <= 114447) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114448 && (row * 640 + col) <= 114559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114560 && (row * 640 + col) <= 114605) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114606 && (row * 640 + col) <= 114625) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114626 && (row * 640 + col) <= 114697) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 114698 && (row * 640 + col) <= 114788) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114789 && (row * 640 + col) <= 114795) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114796 && (row * 640 + col) <= 114808) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114809 && (row * 640 + col) <= 114829) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114830 && (row * 640 + col) <= 114851) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114852 && (row * 640 + col) <= 114866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114867 && (row * 640 + col) <= 114895) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114896 && (row * 640 + col) <= 114906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114907 && (row * 640 + col) <= 114932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114933 && (row * 640 + col) <= 114947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 114948 && (row * 640 + col) <= 114972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 114973 && (row * 640 + col) <= 115041) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115042 && (row * 640 + col) <= 115058) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115059 && (row * 640 + col) <= 115064) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115065 && (row * 640 + col) <= 115087) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115088 && (row * 640 + col) <= 115199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115200 && (row * 640 + col) <= 115245) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115246 && (row * 640 + col) <= 115264) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115265 && (row * 640 + col) <= 115337) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115338 && (row * 640 + col) <= 115428) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115429 && (row * 640 + col) <= 115435) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115436 && (row * 640 + col) <= 115448) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115449 && (row * 640 + col) <= 115469) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115470 && (row * 640 + col) <= 115491) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115492 && (row * 640 + col) <= 115506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115507 && (row * 640 + col) <= 115537) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115538 && (row * 640 + col) <= 115543) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115544 && (row * 640 + col) <= 115572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115573 && (row * 640 + col) <= 115587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115588 && (row * 640 + col) <= 115621) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115622 && (row * 640 + col) <= 115681) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115682 && (row * 640 + col) <= 115698) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115699 && (row * 640 + col) <= 115704) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115705 && (row * 640 + col) <= 115727) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115728 && (row * 640 + col) <= 115839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115840 && (row * 640 + col) <= 115885) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 115886 && (row * 640 + col) <= 115903) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 115904 && (row * 640 + col) <= 115977) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 115978 && (row * 640 + col) <= 116068) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116069 && (row * 640 + col) <= 116075) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116076 && (row * 640 + col) <= 116088) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116089 && (row * 640 + col) <= 116109) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116110 && (row * 640 + col) <= 116131) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116132 && (row * 640 + col) <= 116146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116147 && (row * 640 + col) <= 116177) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116178 && (row * 640 + col) <= 116183) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116184 && (row * 640 + col) <= 116212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116213 && (row * 640 + col) <= 116227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116228 && (row * 640 + col) <= 116261) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116262 && (row * 640 + col) <= 116321) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116322 && (row * 640 + col) <= 116338) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116339 && (row * 640 + col) <= 116344) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116345 && (row * 640 + col) <= 116367) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116368 && (row * 640 + col) <= 116479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116480 && (row * 640 + col) <= 116525) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116526 && (row * 640 + col) <= 116541) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116542 && (row * 640 + col) <= 116617) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 116618 && (row * 640 + col) <= 116708) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116709 && (row * 640 + col) <= 116715) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116716 && (row * 640 + col) <= 116728) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116729 && (row * 640 + col) <= 116749) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116750 && (row * 640 + col) <= 116771) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116772 && (row * 640 + col) <= 116786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116787 && (row * 640 + col) <= 116817) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116818 && (row * 640 + col) <= 116823) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116824 && (row * 640 + col) <= 116852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116853 && (row * 640 + col) <= 116867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116868 && (row * 640 + col) <= 116901) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116902 && (row * 640 + col) <= 116961) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116962 && (row * 640 + col) <= 116978) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 116979 && (row * 640 + col) <= 116984) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 116985 && (row * 640 + col) <= 117007) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117008 && (row * 640 + col) <= 117119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117120 && (row * 640 + col) <= 117165) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117166 && (row * 640 + col) <= 117181) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117182 && (row * 640 + col) <= 117257) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 117258 && (row * 640 + col) <= 117348) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117349 && (row * 640 + col) <= 117355) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117356 && (row * 640 + col) <= 117368) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117369 && (row * 640 + col) <= 117389) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117390 && (row * 640 + col) <= 117411) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117412 && (row * 640 + col) <= 117426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117427 && (row * 640 + col) <= 117457) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117458 && (row * 640 + col) <= 117463) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117464 && (row * 640 + col) <= 117492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117493 && (row * 640 + col) <= 117507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117508 && (row * 640 + col) <= 117541) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117542 && (row * 640 + col) <= 117601) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117602 && (row * 640 + col) <= 117618) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117619 && (row * 640 + col) <= 117624) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117625 && (row * 640 + col) <= 117647) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117648 && (row * 640 + col) <= 117759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117760 && (row * 640 + col) <= 117805) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117806 && (row * 640 + col) <= 117820) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117821 && (row * 640 + col) <= 117897) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 117898 && (row * 640 + col) <= 117988) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 117989 && (row * 640 + col) <= 117995) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 117996 && (row * 640 + col) <= 118008) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118009 && (row * 640 + col) <= 118029) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118030 && (row * 640 + col) <= 118051) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118052 && (row * 640 + col) <= 118066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118067 && (row * 640 + col) <= 118097) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118098 && (row * 640 + col) <= 118103) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118104 && (row * 640 + col) <= 118132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118133 && (row * 640 + col) <= 118147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118148 && (row * 640 + col) <= 118181) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118182 && (row * 640 + col) <= 118241) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118242 && (row * 640 + col) <= 118258) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118259 && (row * 640 + col) <= 118264) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118265 && (row * 640 + col) <= 118287) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118288 && (row * 640 + col) <= 118399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118400 && (row * 640 + col) <= 118445) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118446 && (row * 640 + col) <= 118456) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118457 && (row * 640 + col) <= 118536) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 118537 && (row * 640 + col) <= 118537) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118538 && (row * 640 + col) <= 118628) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118629 && (row * 640 + col) <= 118634) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118635 && (row * 640 + col) <= 118648) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118649 && (row * 640 + col) <= 118669) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118670 && (row * 640 + col) <= 118692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118693 && (row * 640 + col) <= 118706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118707 && (row * 640 + col) <= 118737) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118738 && (row * 640 + col) <= 118743) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118744 && (row * 640 + col) <= 118772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118773 && (row * 640 + col) <= 118787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118788 && (row * 640 + col) <= 118821) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118822 && (row * 640 + col) <= 118881) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118882 && (row * 640 + col) <= 118898) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118899 && (row * 640 + col) <= 118904) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 118905 && (row * 640 + col) <= 118927) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 118928 && (row * 640 + col) <= 119039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119040 && (row * 640 + col) <= 119085) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119086 && (row * 640 + col) <= 119095) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119096 && (row * 640 + col) <= 119175) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119176 && (row * 640 + col) <= 119177) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119178 && (row * 640 + col) <= 119288) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119289 && (row * 640 + col) <= 119309) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119310 && (row * 640 + col) <= 119340) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119341 && (row * 640 + col) <= 119346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119347 && (row * 640 + col) <= 119377) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119378 && (row * 640 + col) <= 119383) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119384 && (row * 640 + col) <= 119412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119413 && (row * 640 + col) <= 119427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119428 && (row * 640 + col) <= 119461) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119462 && (row * 640 + col) <= 119521) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119522 && (row * 640 + col) <= 119567) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119568 && (row * 640 + col) <= 119679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119680 && (row * 640 + col) <= 119725) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119726 && (row * 640 + col) <= 119735) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119736 && (row * 640 + col) <= 119747) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119748 && (row * 640 + col) <= 119750) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119751 && (row * 640 + col) <= 119769) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119770 && (row * 640 + col) <= 119781) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119782 && (row * 640 + col) <= 119801) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 119802 && (row * 640 + col) <= 119817) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119818 && (row * 640 + col) <= 119928) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119929 && (row * 640 + col) <= 119949) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119950 && (row * 640 + col) <= 119980) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 119981 && (row * 640 + col) <= 119986) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 119987 && (row * 640 + col) <= 120017) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120018 && (row * 640 + col) <= 120023) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120024 && (row * 640 + col) <= 120052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120053 && (row * 640 + col) <= 120067) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120068 && (row * 640 + col) <= 120101) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120102 && (row * 640 + col) <= 120161) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120162 && (row * 640 + col) <= 120207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120208 && (row * 640 + col) <= 120319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120320 && (row * 640 + col) <= 120365) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120366 && (row * 640 + col) <= 120375) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120376 && (row * 640 + col) <= 120386) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 120387 && (row * 640 + col) <= 120390) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120391 && (row * 640 + col) <= 120409) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 120410 && (row * 640 + col) <= 120421) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120422 && (row * 640 + col) <= 120441) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 120442 && (row * 640 + col) <= 120457) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120458 && (row * 640 + col) <= 120568) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120569 && (row * 640 + col) <= 120589) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120590 && (row * 640 + col) <= 120620) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120621 && (row * 640 + col) <= 120626) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120627 && (row * 640 + col) <= 120657) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120658 && (row * 640 + col) <= 120663) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120664 && (row * 640 + col) <= 120692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120693 && (row * 640 + col) <= 120707) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120708 && (row * 640 + col) <= 120741) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120742 && (row * 640 + col) <= 120801) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120802 && (row * 640 + col) <= 120847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 120848 && (row * 640 + col) <= 120959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 120960 && (row * 640 + col) <= 121005) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121006 && (row * 640 + col) <= 121018) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121019 && (row * 640 + col) <= 121019) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 121020 && (row * 640 + col) <= 121063) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121064 && (row * 640 + col) <= 121064) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 121065 && (row * 640 + col) <= 121072) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121073 && (row * 640 + col) <= 121073) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 121074 && (row * 640 + col) <= 121097) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121098 && (row * 640 + col) <= 121208) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121209 && (row * 640 + col) <= 121229) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121230 && (row * 640 + col) <= 121260) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121261 && (row * 640 + col) <= 121266) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121267 && (row * 640 + col) <= 121297) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121298 && (row * 640 + col) <= 121303) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121304 && (row * 640 + col) <= 121332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121333 && (row * 640 + col) <= 121347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121348 && (row * 640 + col) <= 121381) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121382 && (row * 640 + col) <= 121441) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121442 && (row * 640 + col) <= 121487) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121488 && (row * 640 + col) <= 121599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121600 && (row * 640 + col) <= 121645) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121646 && (row * 640 + col) <= 121737) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121738 && (row * 640 + col) <= 121848) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121849 && (row * 640 + col) <= 121869) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121870 && (row * 640 + col) <= 121900) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121901 && (row * 640 + col) <= 121906) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121907 && (row * 640 + col) <= 121937) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121938 && (row * 640 + col) <= 121943) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121944 && (row * 640 + col) <= 121972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 121973 && (row * 640 + col) <= 121987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 121988 && (row * 640 + col) <= 122021) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122022 && (row * 640 + col) <= 122081) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122082 && (row * 640 + col) <= 122127) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122128 && (row * 640 + col) <= 122239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122240 && (row * 640 + col) <= 122285) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122286 && (row * 640 + col) <= 122314) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122315 && (row * 640 + col) <= 122318) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122319 && (row * 640 + col) <= 122324) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122325 && (row * 640 + col) <= 122327) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122328 && (row * 640 + col) <= 122341) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122342 && (row * 640 + col) <= 122342) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122343 && (row * 640 + col) <= 122343) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122344 && (row * 640 + col) <= 122344) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122345 && (row * 640 + col) <= 122377) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122378 && (row * 640 + col) <= 122488) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122489 && (row * 640 + col) <= 122509) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122510 && (row * 640 + col) <= 122540) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122541 && (row * 640 + col) <= 122546) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122547 && (row * 640 + col) <= 122577) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122578 && (row * 640 + col) <= 122583) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122584 && (row * 640 + col) <= 122612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122613 && (row * 640 + col) <= 122627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122628 && (row * 640 + col) <= 122661) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122662 && (row * 640 + col) <= 122668) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122669 && (row * 640 + col) <= 122688) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122689 && (row * 640 + col) <= 122689) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122690 && (row * 640 + col) <= 122692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122693 && (row * 640 + col) <= 122703) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122704 && (row * 640 + col) <= 122705) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122706 && (row * 640 + col) <= 122707) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122708 && (row * 640 + col) <= 122709) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122710 && (row * 640 + col) <= 122710) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122711 && (row * 640 + col) <= 122767) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122768 && (row * 640 + col) <= 122879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122880 && (row * 640 + col) <= 122925) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122926 && (row * 640 + col) <= 122954) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 122955 && (row * 640 + col) <= 122985) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 122986 && (row * 640 + col) <= 123017) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123018 && (row * 640 + col) <= 123128) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123129 && (row * 640 + col) <= 123149) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123150 && (row * 640 + col) <= 123180) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123181 && (row * 640 + col) <= 123186) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123187 && (row * 640 + col) <= 123217) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123218 && (row * 640 + col) <= 123223) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123224 && (row * 640 + col) <= 123252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123253 && (row * 640 + col) <= 123267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123268 && (row * 640 + col) <= 123301) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123302 && (row * 640 + col) <= 123307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123308 && (row * 640 + col) <= 123332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123333 && (row * 640 + col) <= 123341) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123342 && (row * 640 + col) <= 123407) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123408 && (row * 640 + col) <= 123519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123520 && (row * 640 + col) <= 123565) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123566 && (row * 640 + col) <= 123594) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123595 && (row * 640 + col) <= 123625) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123626 && (row * 640 + col) <= 123657) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123658 && (row * 640 + col) <= 123768) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123769 && (row * 640 + col) <= 123789) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123790 && (row * 640 + col) <= 123820) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123821 && (row * 640 + col) <= 123826) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123827 && (row * 640 + col) <= 123857) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123858 && (row * 640 + col) <= 123863) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123864 && (row * 640 + col) <= 123892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123893 && (row * 640 + col) <= 123907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123908 && (row * 640 + col) <= 123941) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123942 && (row * 640 + col) <= 123947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123948 && (row * 640 + col) <= 123972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 123973 && (row * 640 + col) <= 123981) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 123982 && (row * 640 + col) <= 124047) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124048 && (row * 640 + col) <= 124159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124160 && (row * 640 + col) <= 124205) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124206 && (row * 640 + col) <= 124234) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124235 && (row * 640 + col) <= 124265) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124266 && (row * 640 + col) <= 124297) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124298 && (row * 640 + col) <= 124409) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124410 && (row * 640 + col) <= 124429) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124430 && (row * 640 + col) <= 124460) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124461 && (row * 640 + col) <= 124466) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124467 && (row * 640 + col) <= 124497) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124498 && (row * 640 + col) <= 124501) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124502 && (row * 640 + col) <= 124502) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124503 && (row * 640 + col) <= 124503) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124504 && (row * 640 + col) <= 124532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124533 && (row * 640 + col) <= 124547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124548 && (row * 640 + col) <= 124581) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124582 && (row * 640 + col) <= 124587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124588 && (row * 640 + col) <= 124612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124613 && (row * 640 + col) <= 124621) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124622 && (row * 640 + col) <= 124687) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124688 && (row * 640 + col) <= 124799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124800 && (row * 640 + col) <= 124845) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124846 && (row * 640 + col) <= 124874) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124875 && (row * 640 + col) <= 124905) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 124906 && (row * 640 + col) <= 124937) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 124938 && (row * 640 + col) <= 125051) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125052 && (row * 640 + col) <= 125069) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125070 && (row * 640 + col) <= 125100) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125101 && (row * 640 + col) <= 125106) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125107 && (row * 640 + col) <= 125137) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125138 && (row * 640 + col) <= 125141) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125142 && (row * 640 + col) <= 125172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125173 && (row * 640 + col) <= 125187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125188 && (row * 640 + col) <= 125221) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125222 && (row * 640 + col) <= 125227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125228 && (row * 640 + col) <= 125252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125253 && (row * 640 + col) <= 125261) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125262 && (row * 640 + col) <= 125327) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125328 && (row * 640 + col) <= 125439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125440 && (row * 640 + col) <= 125485) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125486 && (row * 640 + col) <= 125514) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125515 && (row * 640 + col) <= 125545) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125546 && (row * 640 + col) <= 125577) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125578 && (row * 640 + col) <= 125691) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125692 && (row * 640 + col) <= 125709) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125710 && (row * 640 + col) <= 125740) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125741 && (row * 640 + col) <= 125746) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125747 && (row * 640 + col) <= 125777) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125778 && (row * 640 + col) <= 125781) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125782 && (row * 640 + col) <= 125812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125813 && (row * 640 + col) <= 125827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125828 && (row * 640 + col) <= 125861) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125862 && (row * 640 + col) <= 125867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125868 && (row * 640 + col) <= 125892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125893 && (row * 640 + col) <= 125901) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 125902 && (row * 640 + col) <= 125967) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 125968 && (row * 640 + col) <= 126079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126080 && (row * 640 + col) <= 126125) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126126 && (row * 640 + col) <= 126154) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126155 && (row * 640 + col) <= 126185) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126186 && (row * 640 + col) <= 126217) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126218 && (row * 640 + col) <= 126331) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126332 && (row * 640 + col) <= 126349) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126350 && (row * 640 + col) <= 126380) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126381 && (row * 640 + col) <= 126386) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126387 && (row * 640 + col) <= 126417) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126418 && (row * 640 + col) <= 126421) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126422 && (row * 640 + col) <= 126501) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126502 && (row * 640 + col) <= 126507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126508 && (row * 640 + col) <= 126532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126533 && (row * 640 + col) <= 126541) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126542 && (row * 640 + col) <= 126607) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126608 && (row * 640 + col) <= 126719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126720 && (row * 640 + col) <= 126765) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126766 && (row * 640 + col) <= 126794) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126795 && (row * 640 + col) <= 126825) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126826 && (row * 640 + col) <= 126857) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126858 && (row * 640 + col) <= 126971) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 126972 && (row * 640 + col) <= 126989) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 126990 && (row * 640 + col) <= 127020) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127021 && (row * 640 + col) <= 127026) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127027 && (row * 640 + col) <= 127057) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127058 && (row * 640 + col) <= 127061) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127062 && (row * 640 + col) <= 127141) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127142 && (row * 640 + col) <= 127147) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127148 && (row * 640 + col) <= 127172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127173 && (row * 640 + col) <= 127181) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127182 && (row * 640 + col) <= 127247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127248 && (row * 640 + col) <= 127359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127360 && (row * 640 + col) <= 127405) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127406 && (row * 640 + col) <= 127434) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127435 && (row * 640 + col) <= 127465) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127466 && (row * 640 + col) <= 127497) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127498 && (row * 640 + col) <= 127611) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127612 && (row * 640 + col) <= 127629) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127630 && (row * 640 + col) <= 127660) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127661 && (row * 640 + col) <= 127666) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127667 && (row * 640 + col) <= 127697) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127698 && (row * 640 + col) <= 127701) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127702 && (row * 640 + col) <= 127781) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127782 && (row * 640 + col) <= 127787) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127788 && (row * 640 + col) <= 127812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127813 && (row * 640 + col) <= 127821) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 127822 && (row * 640 + col) <= 127887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 127888 && (row * 640 + col) <= 127999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128000 && (row * 640 + col) <= 128045) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128046 && (row * 640 + col) <= 128071) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128072 && (row * 640 + col) <= 128108) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128109 && (row * 640 + col) <= 128137) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128138 && (row * 640 + col) <= 128251) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128252 && (row * 640 + col) <= 128269) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128270 && (row * 640 + col) <= 128300) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128301 && (row * 640 + col) <= 128306) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128307 && (row * 640 + col) <= 128421) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128422 && (row * 640 + col) <= 128427) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128428 && (row * 640 + col) <= 128452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128453 && (row * 640 + col) <= 128461) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128462 && (row * 640 + col) <= 128527) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128528 && (row * 640 + col) <= 128639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128640 && (row * 640 + col) <= 128685) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128686 && (row * 640 + col) <= 128711) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128712 && (row * 640 + col) <= 128748) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128749 && (row * 640 + col) <= 128777) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128778 && (row * 640 + col) <= 128891) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128892 && (row * 640 + col) <= 128909) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128910 && (row * 640 + col) <= 128940) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 128941 && (row * 640 + col) <= 128946) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 128947 && (row * 640 + col) <= 129061) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129062 && (row * 640 + col) <= 129067) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129068 && (row * 640 + col) <= 129092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129093 && (row * 640 + col) <= 129101) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129102 && (row * 640 + col) <= 129167) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129168 && (row * 640 + col) <= 129279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129280 && (row * 640 + col) <= 129325) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129326 && (row * 640 + col) <= 129351) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129352 && (row * 640 + col) <= 129388) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129389 && (row * 640 + col) <= 129417) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129418 && (row * 640 + col) <= 129531) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129532 && (row * 640 + col) <= 129549) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129550 && (row * 640 + col) <= 129580) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129581 && (row * 640 + col) <= 129586) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129587 && (row * 640 + col) <= 129701) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129702 && (row * 640 + col) <= 129707) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129708 && (row * 640 + col) <= 129732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129733 && (row * 640 + col) <= 129741) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129742 && (row * 640 + col) <= 129807) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129808 && (row * 640 + col) <= 129919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129920 && (row * 640 + col) <= 129965) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 129966 && (row * 640 + col) <= 129991) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 129992 && (row * 640 + col) <= 130028) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130029 && (row * 640 + col) <= 130057) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130058 && (row * 640 + col) <= 130171) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130172 && (row * 640 + col) <= 130180) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130181 && (row * 640 + col) <= 130186) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130187 && (row * 640 + col) <= 130189) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130190 && (row * 640 + col) <= 130223) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130224 && (row * 640 + col) <= 130226) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130227 && (row * 640 + col) <= 130341) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130342 && (row * 640 + col) <= 130347) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130348 && (row * 640 + col) <= 130372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130373 && (row * 640 + col) <= 130381) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130382 && (row * 640 + col) <= 130447) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130448 && (row * 640 + col) <= 130559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130560 && (row * 640 + col) <= 130605) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130606 && (row * 640 + col) <= 130631) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130632 && (row * 640 + col) <= 130668) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130669 && (row * 640 + col) <= 130697) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130698 && (row * 640 + col) <= 130811) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130812 && (row * 640 + col) <= 130820) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130821 && (row * 640 + col) <= 130826) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130827 && (row * 640 + col) <= 130829) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130830 && (row * 640 + col) <= 130863) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130864 && (row * 640 + col) <= 130866) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130867 && (row * 640 + col) <= 130981) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 130982 && (row * 640 + col) <= 130987) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 130988 && (row * 640 + col) <= 131012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131013 && (row * 640 + col) <= 131021) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131022 && (row * 640 + col) <= 131087) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131088 && (row * 640 + col) <= 131199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131200 && (row * 640 + col) <= 131245) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131246 && (row * 640 + col) <= 131271) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131272 && (row * 640 + col) <= 131308) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131309 && (row * 640 + col) <= 131337) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131338 && (row * 640 + col) <= 131451) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131452 && (row * 640 + col) <= 131460) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131461 && (row * 640 + col) <= 131466) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131467 && (row * 640 + col) <= 131469) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131470 && (row * 640 + col) <= 131503) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131504 && (row * 640 + col) <= 131506) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131507 && (row * 640 + col) <= 131621) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131622 && (row * 640 + col) <= 131627) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131628 && (row * 640 + col) <= 131652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131653 && (row * 640 + col) <= 131661) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131662 && (row * 640 + col) <= 131727) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131728 && (row * 640 + col) <= 131839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131840 && (row * 640 + col) <= 131885) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131886 && (row * 640 + col) <= 131911) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131912 && (row * 640 + col) <= 131948) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 131949 && (row * 640 + col) <= 131977) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 131978 && (row * 640 + col) <= 132091) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132092 && (row * 640 + col) <= 132098) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132099 && (row * 640 + col) <= 132143) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132144 && (row * 640 + col) <= 132146) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132147 && (row * 640 + col) <= 132261) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132262 && (row * 640 + col) <= 132267) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132268 && (row * 640 + col) <= 132292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132293 && (row * 640 + col) <= 132301) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132302 && (row * 640 + col) <= 132367) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132368 && (row * 640 + col) <= 132479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132480 && (row * 640 + col) <= 132525) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132526 && (row * 640 + col) <= 132551) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132552 && (row * 640 + col) <= 132588) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132589 && (row * 640 + col) <= 132617) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132618 && (row * 640 + col) <= 132731) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132732 && (row * 640 + col) <= 132737) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132738 && (row * 640 + col) <= 132783) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132784 && (row * 640 + col) <= 132786) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132787 && (row * 640 + col) <= 132901) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132902 && (row * 640 + col) <= 132907) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132908 && (row * 640 + col) <= 132932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 132933 && (row * 640 + col) <= 132941) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 132942 && (row * 640 + col) <= 133007) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133008 && (row * 640 + col) <= 133119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133120 && (row * 640 + col) <= 133165) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133166 && (row * 640 + col) <= 133191) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133192 && (row * 640 + col) <= 133228) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133229 && (row * 640 + col) <= 133257) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133258 && (row * 640 + col) <= 133371) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133372 && (row * 640 + col) <= 133377) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133378 && (row * 640 + col) <= 133423) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133424 && (row * 640 + col) <= 133426) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133427 && (row * 640 + col) <= 133541) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133542 && (row * 640 + col) <= 133547) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133548 && (row * 640 + col) <= 133572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133573 && (row * 640 + col) <= 133581) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133582 && (row * 640 + col) <= 133647) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133648 && (row * 640 + col) <= 133698) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133699 && (row * 640 + col) <= 133708) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 133709 && (row * 640 + col) <= 133759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133760 && (row * 640 + col) <= 133805) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133806 && (row * 640 + col) <= 133831) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133832 && (row * 640 + col) <= 133868) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133869 && (row * 640 + col) <= 133880) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133881 && (row * 640 + col) <= 133888) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 133889 && (row * 640 + col) <= 133897) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 133898 && (row * 640 + col) <= 134063) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134064 && (row * 640 + col) <= 134066) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134067 && (row * 640 + col) <= 134181) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134182 && (row * 640 + col) <= 134187) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134188 && (row * 640 + col) <= 134287) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134288 && (row * 640 + col) <= 134338) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134339 && (row * 640 + col) <= 134349) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 134350 && (row * 640 + col) <= 134399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134400 && (row * 640 + col) <= 134445) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134446 && (row * 640 + col) <= 134471) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134472 && (row * 640 + col) <= 134508) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134509 && (row * 640 + col) <= 134520) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134521 && (row * 640 + col) <= 134528) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134529 && (row * 640 + col) <= 134537) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134538 && (row * 640 + col) <= 134703) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134704 && (row * 640 + col) <= 134706) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134707 && (row * 640 + col) <= 134821) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134822 && (row * 640 + col) <= 134827) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134828 && (row * 640 + col) <= 134927) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 134928 && (row * 640 + col) <= 134977) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134978 && (row * 640 + col) <= 134989) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 134990 && (row * 640 + col) <= 134993) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 134994 && (row * 640 + col) <= 134996) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 134997 && (row * 640 + col) <= 135039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135040 && (row * 640 + col) <= 135085) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135086 && (row * 640 + col) <= 135111) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135112 && (row * 640 + col) <= 135148) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135149 && (row * 640 + col) <= 135159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135160 && (row * 640 + col) <= 135168) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135169 && (row * 640 + col) <= 135177) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135178 && (row * 640 + col) <= 135343) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135344 && (row * 640 + col) <= 135346) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135347 && (row * 640 + col) <= 135461) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135462 && (row * 640 + col) <= 135467) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135468 && (row * 640 + col) <= 135567) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135568 && (row * 640 + col) <= 135615) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135616 && (row * 640 + col) <= 135637) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 135638 && (row * 640 + col) <= 135679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135680 && (row * 640 + col) <= 135725) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135726 && (row * 640 + col) <= 135748) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135749 && (row * 640 + col) <= 135788) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 135789 && (row * 640 + col) <= 135791) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 135792 && (row * 640 + col) <= 136101) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136102 && (row * 640 + col) <= 136107) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136108 && (row * 640 + col) <= 136207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136208 && (row * 640 + col) <= 136222) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136223 && (row * 640 + col) <= 136227) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136228 && (row * 640 + col) <= 136255) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136256 && (row * 640 + col) <= 136277) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 136278 && (row * 640 + col) <= 136319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136320 && (row * 640 + col) <= 136365) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136366 && (row * 640 + col) <= 136388) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136389 && (row * 640 + col) <= 136428) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136429 && (row * 640 + col) <= 136431) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136432 && (row * 640 + col) <= 136741) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136742 && (row * 640 + col) <= 136747) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136748 && (row * 640 + col) <= 136847) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136848 && (row * 640 + col) <= 136862) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136863 && (row * 640 + col) <= 136867) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 136868 && (row * 640 + col) <= 136894) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136895 && (row * 640 + col) <= 136918) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 136919 && (row * 640 + col) <= 136959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 136960 && (row * 640 + col) <= 137005) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 137006 && (row * 640 + col) <= 137028) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137029 && (row * 640 + col) <= 137068) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 137069 && (row * 640 + col) <= 137071) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137072 && (row * 640 + col) <= 137381) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 137382 && (row * 640 + col) <= 137387) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137388 && (row * 640 + col) <= 137487) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 137488 && (row * 640 + col) <= 137501) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137502 && (row * 640 + col) <= 137508) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 137509 && (row * 640 + col) <= 137532) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137533 && (row * 640 + col) <= 137560) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 137561 && (row * 640 + col) <= 137599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137600 && (row * 640 + col) <= 137645) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 137646 && (row * 640 + col) <= 137668) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137669 && (row * 640 + col) <= 137708) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 137709 && (row * 640 + col) <= 137711) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 137712 && (row * 640 + col) <= 138021) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138022 && (row * 640 + col) <= 138027) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138028 && (row * 640 + col) <= 138156) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138157 && (row * 640 + col) <= 138172) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138173 && (row * 640 + col) <= 138200) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 138201 && (row * 640 + col) <= 138239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138240 && (row * 640 + col) <= 138285) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138286 && (row * 640 + col) <= 138308) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138309 && (row * 640 + col) <= 138348) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138349 && (row * 640 + col) <= 138351) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138352 && (row * 640 + col) <= 138661) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138662 && (row * 640 + col) <= 138667) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138668 && (row * 640 + col) <= 138796) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138797 && (row * 640 + col) <= 138799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138800 && (row * 640 + col) <= 138840) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 138841 && (row * 640 + col) <= 138879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138880 && (row * 640 + col) <= 138925) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138926 && (row * 640 + col) <= 138948) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138949 && (row * 640 + col) <= 138988) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 138989 && (row * 640 + col) <= 138991) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 138992 && (row * 640 + col) <= 139301) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 139302 && (row * 640 + col) <= 139307) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 139308 && (row * 640 + col) <= 139436) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 139437 && (row * 640 + col) <= 139438) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 139439 && (row * 640 + col) <= 139480) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 139481 && (row * 640 + col) <= 139519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 139520 && (row * 640 + col) <= 139565) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 139566 && (row * 640 + col) <= 139588) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 139589 && (row * 640 + col) <= 139628) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 139629 && (row * 640 + col) <= 139631) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 139632 && (row * 640 + col) <= 139941) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 139942 && (row * 640 + col) <= 139947) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 139948 && (row * 640 + col) <= 140076) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 140077 && (row * 640 + col) <= 140078) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140079 && (row * 640 + col) <= 140120) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 140121 && (row * 640 + col) <= 140159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140160 && (row * 640 + col) <= 140205) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 140206 && (row * 640 + col) <= 140228) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140229 && (row * 640 + col) <= 140268) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 140269 && (row * 640 + col) <= 140271) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140272 && (row * 640 + col) <= 140581) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 140582 && (row * 640 + col) <= 140587) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140588 && (row * 640 + col) <= 140716) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 140717 && (row * 640 + col) <= 140764) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 140765 && (row * 640 + col) <= 140799) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140800 && (row * 640 + col) <= 140850) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 140851 && (row * 640 + col) <= 140859) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140860 && (row * 640 + col) <= 140908) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 140909 && (row * 640 + col) <= 140911) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 140912 && (row * 640 + col) <= 141221) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 141222 && (row * 640 + col) <= 141227) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 141228 && (row * 640 + col) <= 141356) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 141357 && (row * 640 + col) <= 141405) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 141406 && (row * 640 + col) <= 141439) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 141440 && (row * 640 + col) <= 141490) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 141491 && (row * 640 + col) <= 141499) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 141500 && (row * 640 + col) <= 141548) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 141549 && (row * 640 + col) <= 141551) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 141552 && (row * 640 + col) <= 141861) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 141862 && (row * 640 + col) <= 141867) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 141868 && (row * 640 + col) <= 141996) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 141997 && (row * 640 + col) <= 142046) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 142047 && (row * 640 + col) <= 142079) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 142080 && (row * 640 + col) <= 142130) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 142131 && (row * 640 + col) <= 142139) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 142140 && (row * 640 + col) <= 142188) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 142189 && (row * 640 + col) <= 142191) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 142192 && (row * 640 + col) <= 142501) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 142502 && (row * 640 + col) <= 142507) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 142508 && (row * 640 + col) <= 142636) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 142637 && (row * 640 + col) <= 142690) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 142691 && (row * 640 + col) <= 142719) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 142720 && (row * 640 + col) <= 142770) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 142771 && (row * 640 + col) <= 142779) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 142780 && (row * 640 + col) <= 142828) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 142829 && (row * 640 + col) <= 142831) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 142832 && (row * 640 + col) <= 143276) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 143277 && (row * 640 + col) <= 143331) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 143332 && (row * 640 + col) <= 143359) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 143360 && (row * 640 + col) <= 143410) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 143411 && (row * 640 + col) <= 143419) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 143420 && (row * 640 + col) <= 143468) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 143469 && (row * 640 + col) <= 143471) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 143472 && (row * 640 + col) <= 143916) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 143917 && (row * 640 + col) <= 143971) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 143972 && (row * 640 + col) <= 143999) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 144000 && (row * 640 + col) <= 144050) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 144051 && (row * 640 + col) <= 144059) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 144060 && (row * 640 + col) <= 144108) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 144109 && (row * 640 + col) <= 144111) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 144112 && (row * 640 + col) <= 144556) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 144557 && (row * 640 + col) <= 144611) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 144612 && (row * 640 + col) <= 144639) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 144640 && (row * 640 + col) <= 144690) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 144691 && (row * 640 + col) <= 144699) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 144700 && (row * 640 + col) <= 144748) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 144749 && (row * 640 + col) <= 144751) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 144752 && (row * 640 + col) <= 145196) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 145197 && (row * 640 + col) <= 145197) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145198 && (row * 640 + col) <= 145250) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 145251 && (row * 640 + col) <= 145279) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145280 && (row * 640 + col) <= 145330) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 145331 && (row * 640 + col) <= 145339) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145340 && (row * 640 + col) <= 145388) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 145389 && (row * 640 + col) <= 145391) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145392 && (row * 640 + col) <= 145836) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 145837 && (row * 640 + col) <= 145919) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145920 && (row * 640 + col) <= 145970) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 145971 && (row * 640 + col) <= 145979) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 145980 && (row * 640 + col) <= 146028) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 146029 && (row * 640 + col) <= 146031) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 146032 && (row * 640 + col) <= 146476) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 146477 && (row * 640 + col) <= 146559) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 146560 && (row * 640 + col) <= 146610) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 146611 && (row * 640 + col) <= 146619) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 146620 && (row * 640 + col) <= 147116) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 147117 && (row * 640 + col) <= 147199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 147200 && (row * 640 + col) <= 147250) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 147251 && (row * 640 + col) <= 147259) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 147260 && (row * 640 + col) <= 147478) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 147479 && (row * 640 + col) <= 147483) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 147484 && (row * 640 + col) <= 147756) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 147757 && (row * 640 + col) <= 147839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 147840 && (row * 640 + col) <= 147891) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 147892 && (row * 640 + col) <= 147899) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 147900 && (row * 640 + col) <= 148118) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 148119 && (row * 640 + col) <= 148147) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 148148 && (row * 640 + col) <= 148396) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 148397 && (row * 640 + col) <= 148479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 148480 && (row * 640 + col) <= 148692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 148693 && (row * 640 + col) <= 148695) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 148696 && (row * 640 + col) <= 148758) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 148759 && (row * 640 + col) <= 148789) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 148790 && (row * 640 + col) <= 149036) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149037 && (row * 640 + col) <= 149085) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149086 && (row * 640 + col) <= 149087) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149088 && (row * 640 + col) <= 149119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149120 && (row * 640 + col) <= 149332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149333 && (row * 640 + col) <= 149335) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 149336 && (row * 640 + col) <= 149398) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149399 && (row * 640 + col) <= 149431) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 149432 && (row * 640 + col) <= 149676) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149677 && (row * 640 + col) <= 149725) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149726 && (row * 640 + col) <= 149727) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149728 && (row * 640 + col) <= 149759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 149760 && (row * 640 + col) <= 149972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 149973 && (row * 640 + col) <= 149975) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 149976 && (row * 640 + col) <= 150038) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150039 && (row * 640 + col) <= 150041) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 150042 && (row * 640 + col) <= 150064) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150065 && (row * 640 + col) <= 150072) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 150073 && (row * 640 + col) <= 150316) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150317 && (row * 640 + col) <= 150364) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 150365 && (row * 640 + col) <= 150368) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150369 && (row * 640 + col) <= 150399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 150400 && (row * 640 + col) <= 150612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150613 && (row * 640 + col) <= 150615) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 150616 && (row * 640 + col) <= 150678) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150679 && (row * 640 + col) <= 150681) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 150682 && (row * 640 + col) <= 150707) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150708 && (row * 640 + col) <= 150713) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 150714 && (row * 640 + col) <= 150956) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 150957 && (row * 640 + col) <= 151002) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151003 && (row * 640 + col) <= 151010) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151011 && (row * 640 + col) <= 151033) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151034 && (row * 640 + col) <= 151034) color_data <= 12'b000001111110; else
        if ((row * 640 + col) >= 151035 && (row * 640 + col) <= 151252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151253 && (row * 640 + col) <= 151255) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151256 && (row * 640 + col) <= 151318) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151319 && (row * 640 + col) <= 151321) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151322 && (row * 640 + col) <= 151348) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151349 && (row * 640 + col) <= 151353) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151354 && (row * 640 + col) <= 151596) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151597 && (row * 640 + col) <= 151642) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151643 && (row * 640 + col) <= 151650) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151651 && (row * 640 + col) <= 151673) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 151674 && (row * 640 + col) <= 151674) color_data <= 12'b000001111110; else
        if ((row * 640 + col) >= 151675 && (row * 640 + col) <= 151892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151893 && (row * 640 + col) <= 151895) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151896 && (row * 640 + col) <= 151958) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151959 && (row * 640 + col) <= 151961) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151962 && (row * 640 + col) <= 151989) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 151990 && (row * 640 + col) <= 151993) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 151994 && (row * 640 + col) <= 152236) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152237 && (row * 640 + col) <= 152282) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152283 && (row * 640 + col) <= 152290) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152291 && (row * 640 + col) <= 152313) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152314 && (row * 640 + col) <= 152314) color_data <= 12'b000001111110; else
        if ((row * 640 + col) >= 152315 && (row * 640 + col) <= 152532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152533 && (row * 640 + col) <= 152535) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 152536 && (row * 640 + col) <= 152598) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152599 && (row * 640 + col) <= 152601) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 152602 && (row * 640 + col) <= 152630) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152631 && (row * 640 + col) <= 152633) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 152634 && (row * 640 + col) <= 152876) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152877 && (row * 640 + col) <= 152899) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152900 && (row * 640 + col) <= 152904) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152905 && (row * 640 + col) <= 152922) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152923 && (row * 640 + col) <= 152930) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 152931 && (row * 640 + col) <= 152953) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 152954 && (row * 640 + col) <= 152954) color_data <= 12'b000001111110; else
        if ((row * 640 + col) >= 152955 && (row * 640 + col) <= 153172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153173 && (row * 640 + col) <= 153175) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 153176 && (row * 640 + col) <= 153238) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153239 && (row * 640 + col) <= 153241) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 153242 && (row * 640 + col) <= 153270) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153271 && (row * 640 + col) <= 153273) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 153274 && (row * 640 + col) <= 153516) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153517 && (row * 640 + col) <= 153539) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153540 && (row * 640 + col) <= 153544) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153545 && (row * 640 + col) <= 153562) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153563 && (row * 640 + col) <= 153570) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153571 && (row * 640 + col) <= 153593) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 153594 && (row * 640 + col) <= 153594) color_data <= 12'b000001111110; else
        if ((row * 640 + col) >= 153595 && (row * 640 + col) <= 153812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153813 && (row * 640 + col) <= 153815) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 153816 && (row * 640 + col) <= 153878) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153879 && (row * 640 + col) <= 153881) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 153882 && (row * 640 + col) <= 153909) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 153910 && (row * 640 + col) <= 153913) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 153914 && (row * 640 + col) <= 154156) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154157 && (row * 640 + col) <= 154179) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154180 && (row * 640 + col) <= 154184) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154185 && (row * 640 + col) <= 154199) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154200 && (row * 640 + col) <= 154452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154453 && (row * 640 + col) <= 154455) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 154456 && (row * 640 + col) <= 154495) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154496 && (row * 640 + col) <= 154498) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 154499 && (row * 640 + col) <= 154518) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154519 && (row * 640 + col) <= 154521) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 154522 && (row * 640 + col) <= 154548) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154549 && (row * 640 + col) <= 154553) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 154554 && (row * 640 + col) <= 154796) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154797 && (row * 640 + col) <= 154819) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154820 && (row * 640 + col) <= 154824) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 154825 && (row * 640 + col) <= 154839) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 154840 && (row * 640 + col) <= 155092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155093 && (row * 640 + col) <= 155095) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155096 && (row * 640 + col) <= 155135) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155136 && (row * 640 + col) <= 155138) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155139 && (row * 640 + col) <= 155158) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155159 && (row * 640 + col) <= 155161) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155162 && (row * 640 + col) <= 155186) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155187 && (row * 640 + col) <= 155193) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155194 && (row * 640 + col) <= 155436) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155437 && (row * 640 + col) <= 155459) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155460 && (row * 640 + col) <= 155464) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155465 && (row * 640 + col) <= 155479) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 155480 && (row * 640 + col) <= 155732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155733 && (row * 640 + col) <= 155735) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155736 && (row * 640 + col) <= 155775) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155776 && (row * 640 + col) <= 155778) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155779 && (row * 640 + col) <= 155798) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155799 && (row * 640 + col) <= 155801) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155802 && (row * 640 + col) <= 155825) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 155826 && (row * 640 + col) <= 155832) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 155833 && (row * 640 + col) <= 156076) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156077 && (row * 640 + col) <= 156087) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156088 && (row * 640 + col) <= 156110) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156111 && (row * 640 + col) <= 156119) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156120 && (row * 640 + col) <= 156372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156373 && (row * 640 + col) <= 156375) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 156376 && (row * 640 + col) <= 156415) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156416 && (row * 640 + col) <= 156418) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 156419 && (row * 640 + col) <= 156438) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156439 && (row * 640 + col) <= 156441) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 156442 && (row * 640 + col) <= 156462) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156463 && (row * 640 + col) <= 156471) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 156472 && (row * 640 + col) <= 156716) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156717 && (row * 640 + col) <= 156727) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156728 && (row * 640 + col) <= 156750) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 156751 && (row * 640 + col) <= 156759) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 156760 && (row * 640 + col) <= 157012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157013 && (row * 640 + col) <= 157015) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157016 && (row * 640 + col) <= 157055) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157056 && (row * 640 + col) <= 157058) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157059 && (row * 640 + col) <= 157078) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157079 && (row * 640 + col) <= 157081) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157082 && (row * 640 + col) <= 157098) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157099 && (row * 640 + col) <= 157109) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157110 && (row * 640 + col) <= 157356) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157357 && (row * 640 + col) <= 157367) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157368 && (row * 640 + col) <= 157390) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157391 && (row * 640 + col) <= 157399) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 157400 && (row * 640 + col) <= 157652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157653 && (row * 640 + col) <= 157655) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157656 && (row * 640 + col) <= 157695) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157696 && (row * 640 + col) <= 157698) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157699 && (row * 640 + col) <= 157718) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157719 && (row * 640 + col) <= 157721) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157722 && (row * 640 + col) <= 157730) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157731 && (row * 640 + col) <= 157747) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 157748 && (row * 640 + col) <= 157996) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 157997 && (row * 640 + col) <= 158007) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158008 && (row * 640 + col) <= 158030) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158031 && (row * 640 + col) <= 158039) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158040 && (row * 640 + col) <= 158292) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158293 && (row * 640 + col) <= 158295) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 158296 && (row * 640 + col) <= 158335) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158336 && (row * 640 + col) <= 158338) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 158339 && (row * 640 + col) <= 158358) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158359 && (row * 640 + col) <= 158384) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 158385 && (row * 640 + col) <= 158636) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158637 && (row * 640 + col) <= 158647) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158648 && (row * 640 + col) <= 158670) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158671 && (row * 640 + col) <= 158679) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 158680 && (row * 640 + col) <= 158932) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158933 && (row * 640 + col) <= 158935) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 158936 && (row * 640 + col) <= 158975) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158976 && (row * 640 + col) <= 158978) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 158979 && (row * 640 + col) <= 158998) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 158999 && (row * 640 + col) <= 159020) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 159021 && (row * 640 + col) <= 159276) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159277 && (row * 640 + col) <= 159287) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159288 && (row * 640 + col) <= 159310) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159311 && (row * 640 + col) <= 159319) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159320 && (row * 640 + col) <= 159572) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159573 && (row * 640 + col) <= 159575) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 159576 && (row * 640 + col) <= 159607) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159608 && (row * 640 + col) <= 159627) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 159628 && (row * 640 + col) <= 159638) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159639 && (row * 640 + col) <= 159652) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 159653 && (row * 640 + col) <= 159950) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 159951 && (row * 640 + col) <= 159959) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 159960 && (row * 640 + col) <= 160212) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160213 && (row * 640 + col) <= 160215) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160216 && (row * 640 + col) <= 160247) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160248 && (row * 640 + col) <= 160267) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160268 && (row * 640 + col) <= 160278) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160279 && (row * 640 + col) <= 160288) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160289 && (row * 640 + col) <= 160590) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160591 && (row * 640 + col) <= 160599) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 160600 && (row * 640 + col) <= 160852) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160853 && (row * 640 + col) <= 160855) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160856 && (row * 640 + col) <= 160887) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160888 && (row * 640 + col) <= 160907) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160908 && (row * 640 + col) <= 160918) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160919 && (row * 640 + col) <= 160921) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160922 && (row * 640 + col) <= 160922) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 160923 && (row * 640 + col) <= 160930) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 160931 && (row * 640 + col) <= 161230) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161231 && (row * 640 + col) <= 161239) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161240 && (row * 640 + col) <= 161492) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161493 && (row * 640 + col) <= 161495) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 161496 && (row * 640 + col) <= 161535) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161536 && (row * 640 + col) <= 161538) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 161539 && (row * 640 + col) <= 161558) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161559 && (row * 640 + col) <= 161561) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 161562 && (row * 640 + col) <= 161564) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161565 && (row * 640 + col) <= 161572) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 161573 && (row * 640 + col) <= 161870) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 161871 && (row * 640 + col) <= 161879) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 161880 && (row * 640 + col) <= 162132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162133 && (row * 640 + col) <= 162135) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162136 && (row * 640 + col) <= 162175) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162176 && (row * 640 + col) <= 162178) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162179 && (row * 640 + col) <= 162198) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162199 && (row * 640 + col) <= 162201) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162202 && (row * 640 + col) <= 162207) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162208 && (row * 640 + col) <= 162214) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162215 && (row * 640 + col) <= 162510) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162511 && (row * 640 + col) <= 162519) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 162520 && (row * 640 + col) <= 162772) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162773 && (row * 640 + col) <= 162775) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162776 && (row * 640 + col) <= 162815) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162816 && (row * 640 + col) <= 162818) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162819 && (row * 640 + col) <= 162838) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162839 && (row * 640 + col) <= 162841) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162842 && (row * 640 + col) <= 162848) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 162849 && (row * 640 + col) <= 162855) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 162856 && (row * 640 + col) <= 163150) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 163151 && (row * 640 + col) <= 163159) color_data <= 12'b000110111111; else
        if ((row * 640 + col) >= 163160 && (row * 640 + col) <= 163412) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 163413 && (row * 640 + col) <= 163415) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 163416 && (row * 640 + col) <= 163455) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 163456 && (row * 640 + col) <= 163458) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 163459 && (row * 640 + col) <= 163478) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 163479 && (row * 640 + col) <= 163481) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 163482 && (row * 640 + col) <= 163490) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 163491 && (row * 640 + col) <= 163496) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 163497 && (row * 640 + col) <= 164052) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164053 && (row * 640 + col) <= 164055) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164056 && (row * 640 + col) <= 164095) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164096 && (row * 640 + col) <= 164098) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164099 && (row * 640 + col) <= 164118) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164119 && (row * 640 + col) <= 164121) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164122 && (row * 640 + col) <= 164132) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164133 && (row * 640 + col) <= 164138) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164139 && (row * 640 + col) <= 164692) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164693 && (row * 640 + col) <= 164695) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164696 && (row * 640 + col) <= 164735) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164736 && (row * 640 + col) <= 164738) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164739 && (row * 640 + col) <= 164758) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164759 && (row * 640 + col) <= 164761) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164762 && (row * 640 + col) <= 164773) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 164774 && (row * 640 + col) <= 164780) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 164781 && (row * 640 + col) <= 165332) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 165333 && (row * 640 + col) <= 165335) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165336 && (row * 640 + col) <= 165375) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 165376 && (row * 640 + col) <= 165378) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165379 && (row * 640 + col) <= 165398) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 165399 && (row * 640 + col) <= 165401) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165402 && (row * 640 + col) <= 165415) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 165416 && (row * 640 + col) <= 165421) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165422 && (row * 640 + col) <= 165972) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 165973 && (row * 640 + col) <= 165975) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 165976 && (row * 640 + col) <= 166015) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166016 && (row * 640 + col) <= 166018) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166019 && (row * 640 + col) <= 166038) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166039 && (row * 640 + col) <= 166041) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166042 && (row * 640 + col) <= 166057) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166058 && (row * 640 + col) <= 166062) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166063 && (row * 640 + col) <= 166612) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166613 && (row * 640 + col) <= 166615) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166616 && (row * 640 + col) <= 166655) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166656 && (row * 640 + col) <= 166658) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166659 && (row * 640 + col) <= 166678) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166679 && (row * 640 + col) <= 166681) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166682 && (row * 640 + col) <= 166698) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 166699 && (row * 640 + col) <= 166703) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 166704 && (row * 640 + col) <= 167252) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167253 && (row * 640 + col) <= 167255) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167256 && (row * 640 + col) <= 167295) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167296 && (row * 640 + col) <= 167298) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167299 && (row * 640 + col) <= 167318) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167319 && (row * 640 + col) <= 167321) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167322 && (row * 640 + col) <= 167338) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167339 && (row * 640 + col) <= 167344) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167345 && (row * 640 + col) <= 167892) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167893 && (row * 640 + col) <= 167895) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167896 && (row * 640 + col) <= 167935) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167936 && (row * 640 + col) <= 167938) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167939 && (row * 640 + col) <= 167958) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167959 && (row * 640 + col) <= 167961) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167962 && (row * 640 + col) <= 167980) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 167981 && (row * 640 + col) <= 167985) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 167986 && (row * 640 + col) <= 168532) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 168533 && (row * 640 + col) <= 168535) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 168536 && (row * 640 + col) <= 168598) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 168599 && (row * 640 + col) <= 168601) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 168602 && (row * 640 + col) <= 168621) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 168622 && (row * 640 + col) <= 168626) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 168627 && (row * 640 + col) <= 169172) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 169173 && (row * 640 + col) <= 169175) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 169176 && (row * 640 + col) <= 169238) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 169239 && (row * 640 + col) <= 169241) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 169242 && (row * 640 + col) <= 169262) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 169263 && (row * 640 + col) <= 169267) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 169268 && (row * 640 + col) <= 169812) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 169813 && (row * 640 + col) <= 169815) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 169816 && (row * 640 + col) <= 169878) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 169879 && (row * 640 + col) <= 169881) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 169882 && (row * 640 + col) <= 169903) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 169904 && (row * 640 + col) <= 169907) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 169908 && (row * 640 + col) <= 170452) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 170453 && (row * 640 + col) <= 170455) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 170456 && (row * 640 + col) <= 170518) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 170519 && (row * 640 + col) <= 170521) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 170522 && (row * 640 + col) <= 170543) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 170544 && (row * 640 + col) <= 170548) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 170549 && (row * 640 + col) <= 171092) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171093 && (row * 640 + col) <= 171095) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 171096 && (row * 640 + col) <= 171158) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171159 && (row * 640 + col) <= 171161) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 171162 && (row * 640 + col) <= 171184) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171185 && (row * 640 + col) <= 171189) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 171190 && (row * 640 + col) <= 171732) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171733 && (row * 640 + col) <= 171735) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 171736 && (row * 640 + col) <= 171798) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171799 && (row * 640 + col) <= 171801) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 171802 && (row * 640 + col) <= 171825) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 171826 && (row * 640 + col) <= 171829) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 171830 && (row * 640 + col) <= 172372) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 172373 && (row * 640 + col) <= 172394) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 172395 && (row * 640 + col) <= 172438) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 172439 && (row * 640 + col) <= 172441) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 172442 && (row * 640 + col) <= 172465) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 172466 && (row * 640 + col) <= 172470) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 172471 && (row * 640 + col) <= 173012) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173013 && (row * 640 + col) <= 173034) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173035 && (row * 640 + col) <= 173078) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173079 && (row * 640 + col) <= 173081) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173082 && (row * 640 + col) <= 173106) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173107 && (row * 640 + col) <= 173110) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173111 && (row * 640 + col) <= 173652) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173653 && (row * 640 + col) <= 173674) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173675 && (row * 640 + col) <= 173718) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173719 && (row * 640 + col) <= 173721) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173722 && (row * 640 + col) <= 173747) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 173748 && (row * 640 + col) <= 173751) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 173752 && (row * 640 + col) <= 174358) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 174359 && (row * 640 + col) <= 174361) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 174362 && (row * 640 + col) <= 174387) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 174388 && (row * 640 + col) <= 174391) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 174392 && (row * 640 + col) <= 175028) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 175029 && (row * 640 + col) <= 175031) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 175032 && (row * 640 + col) <= 181119) color_data <= 12'b000001111101; else
        if ((row * 640 + col) >= 181120 && (row * 640 + col) <= 204799) color_data <= 12'b010010000001; else
        if ((row * 640 + col) >= 204800 && (row * 640 + col) <= 207251) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 207252 && (row * 640 + col) <= 207275) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207276 && (row * 640 + col) <= 207887) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 207888 && (row * 640 + col) <= 207917) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 207918 && (row * 640 + col) <= 208520) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 208521 && (row * 640 + col) <= 208562) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 208563 && (row * 640 + col) <= 209154) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 209155 && (row * 640 + col) <= 209207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209208 && (row * 640 + col) <= 209792) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 209793 && (row * 640 + col) <= 209809) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209810 && (row * 640 + col) <= 209812) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 209813 && (row * 640 + col) <= 209848) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 209849 && (row * 640 + col) <= 210273) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 210274 && (row * 640 + col) <= 210279) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210280 && (row * 640 + col) <= 210430) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 210431 && (row * 640 + col) <= 210444) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210445 && (row * 640 + col) <= 210454) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 210455 && (row * 640 + col) <= 210457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210458 && (row * 640 + col) <= 210474) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 210475 && (row * 640 + col) <= 210489) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210490 && (row * 640 + col) <= 210910) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 210911 && (row * 640 + col) <= 210913) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210914 && (row * 640 + col) <= 210919) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 210920 && (row * 640 + col) <= 210922) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 210923 && (row * 640 + col) <= 211069) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 211070 && (row * 640 + col) <= 211082) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211083 && (row * 640 + col) <= 211094) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 211095 && (row * 640 + col) <= 211097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211098 && (row * 640 + col) <= 211118) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 211119 && (row * 640 + col) <= 211130) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211131 && (row * 640 + col) <= 211549) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 211550 && (row * 640 + col) <= 211550) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211551 && (row * 640 + col) <= 211562) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 211563 && (row * 640 + col) <= 211563) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211564 && (row * 640 + col) <= 211708) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 211709 && (row * 640 + col) <= 211718) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211719 && (row * 640 + col) <= 211734) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 211735 && (row * 640 + col) <= 211737) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211738 && (row * 640 + col) <= 211763) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 211764 && (row * 640 + col) <= 211771) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 211772 && (row * 640 + col) <= 212187) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 212188 && (row * 640 + col) <= 212189) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212190 && (row * 640 + col) <= 212203) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 212204 && (row * 640 + col) <= 212205) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212206 && (row * 640 + col) <= 212347) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 212348 && (row * 640 + col) <= 212356) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212357 && (row * 640 + col) <= 212374) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 212375 && (row * 640 + col) <= 212377) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212378 && (row * 640 + col) <= 212405) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 212406 && (row * 640 + col) <= 212411) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212412 && (row * 640 + col) <= 212826) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 212827 && (row * 640 + col) <= 212827) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212828 && (row * 640 + col) <= 212830) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 212831 && (row * 640 + col) <= 212831) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212832 && (row * 640 + col) <= 212834) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 212835 && (row * 640 + col) <= 212835) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212836 && (row * 640 + col) <= 212838) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 212839 && (row * 640 + col) <= 212839) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212840 && (row * 640 + col) <= 212842) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 212843 && (row * 640 + col) <= 212843) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212844 && (row * 640 + col) <= 212845) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 212846 && (row * 640 + col) <= 212846) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212847 && (row * 640 + col) <= 212985) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 212986 && (row * 640 + col) <= 212993) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 212994 && (row * 640 + col) <= 213014) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 213015 && (row * 640 + col) <= 213017) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213018 && (row * 640 + col) <= 213046) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 213047 && (row * 640 + col) <= 213052) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213053 && (row * 640 + col) <= 213466) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 213467 && (row * 640 + col) <= 213467) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213468 && (row * 640 + col) <= 213471) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 213472 && (row * 640 + col) <= 213472) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213473 && (row * 640 + col) <= 213473) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 213474 && (row * 640 + col) <= 213474) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213475 && (row * 640 + col) <= 213479) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 213480 && (row * 640 + col) <= 213480) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213481 && (row * 640 + col) <= 213481) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 213482 && (row * 640 + col) <= 213482) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213483 && (row * 640 + col) <= 213485) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 213486 && (row * 640 + col) <= 213486) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213487 && (row * 640 + col) <= 213624) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 213625 && (row * 640 + col) <= 213631) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213632 && (row * 640 + col) <= 213654) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 213655 && (row * 640 + col) <= 213657) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213658 && (row * 640 + col) <= 213686) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 213687 && (row * 640 + col) <= 213692) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 213693 && (row * 640 + col) <= 214105) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 214106 && (row * 640 + col) <= 214106) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214107 && (row * 640 + col) <= 214112) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214113 && (row * 640 + col) <= 214113) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214114 && (row * 640 + col) <= 214120) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214121 && (row * 640 + col) <= 214121) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214122 && (row * 640 + col) <= 214126) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214127 && (row * 640 + col) <= 214128) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214129 && (row * 640 + col) <= 214263) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 214264 && (row * 640 + col) <= 214270) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214271 && (row * 640 + col) <= 214294) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 214295 && (row * 640 + col) <= 214297) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214298 && (row * 640 + col) <= 214327) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 214328 && (row * 640 + col) <= 214332) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214333 && (row * 640 + col) <= 214745) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 214746 && (row * 640 + col) <= 214746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214747 && (row * 640 + col) <= 214751) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214752 && (row * 640 + col) <= 214752) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214753 && (row * 640 + col) <= 214753) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214754 && (row * 640 + col) <= 214754) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214755 && (row * 640 + col) <= 214759) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214760 && (row * 640 + col) <= 214760) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214761 && (row * 640 + col) <= 214761) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214762 && (row * 640 + col) <= 214762) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214763 && (row * 640 + col) <= 214767) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 214768 && (row * 640 + col) <= 214768) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214769 && (row * 640 + col) <= 214903) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 214904 && (row * 640 + col) <= 214909) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214910 && (row * 640 + col) <= 214934) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 214935 && (row * 640 + col) <= 214937) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214938 && (row * 640 + col) <= 214967) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 214968 && (row * 640 + col) <= 214972) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 214973 && (row * 640 + col) <= 215384) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 215385 && (row * 640 + col) <= 215385) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215386 && (row * 640 + col) <= 215390) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 215391 && (row * 640 + col) <= 215391) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215392 && (row * 640 + col) <= 215394) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 215395 && (row * 640 + col) <= 215395) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215396 && (row * 640 + col) <= 215398) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 215399 && (row * 640 + col) <= 215399) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215400 && (row * 640 + col) <= 215402) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 215403 && (row * 640 + col) <= 215403) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215404 && (row * 640 + col) <= 215407) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 215408 && (row * 640 + col) <= 215408) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215409 && (row * 640 + col) <= 215542) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 215543 && (row * 640 + col) <= 215547) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215548 && (row * 640 + col) <= 215574) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 215575 && (row * 640 + col) <= 215577) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215578 && (row * 640 + col) <= 215608) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 215609 && (row * 640 + col) <= 215612) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 215613 && (row * 640 + col) <= 216024) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 216025 && (row * 640 + col) <= 216025) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216026 && (row * 640 + col) <= 216047) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 216048 && (row * 640 + col) <= 216048) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216049 && (row * 640 + col) <= 216182) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 216183 && (row * 640 + col) <= 216186) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216187 && (row * 640 + col) <= 216214) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 216215 && (row * 640 + col) <= 216217) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216218 && (row * 640 + col) <= 216248) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 216249 && (row * 640 + col) <= 216252) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216253 && (row * 640 + col) <= 216663) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 216664 && (row * 640 + col) <= 216664) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216665 && (row * 640 + col) <= 216688) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 216689 && (row * 640 + col) <= 216689) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216690 && (row * 640 + col) <= 216822) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 216823 && (row * 640 + col) <= 216826) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216827 && (row * 640 + col) <= 216854) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 216855 && (row * 640 + col) <= 216857) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216858 && (row * 640 + col) <= 216888) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 216889 && (row * 640 + col) <= 216893) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 216894 && (row * 640 + col) <= 217303) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 217304 && (row * 640 + col) <= 217304) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217305 && (row * 640 + col) <= 217328) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 217329 && (row * 640 + col) <= 217329) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217330 && (row * 640 + col) <= 217462) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 217463 && (row * 640 + col) <= 217466) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217467 && (row * 640 + col) <= 217494) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 217495 && (row * 640 + col) <= 217497) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217498 && (row * 640 + col) <= 217528) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 217529 && (row * 640 + col) <= 217536) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217537 && (row * 640 + col) <= 217943) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 217944 && (row * 640 + col) <= 217944) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217945 && (row * 640 + col) <= 217968) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 217969 && (row * 640 + col) <= 217969) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 217970 && (row * 640 + col) <= 218102) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 218103 && (row * 640 + col) <= 218106) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218107 && (row * 640 + col) <= 218134) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 218135 && (row * 640 + col) <= 218137) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218138 && (row * 640 + col) <= 218168) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 218169 && (row * 640 + col) <= 218177) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218178 && (row * 640 + col) <= 218583) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 218584 && (row * 640 + col) <= 218584) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218585 && (row * 640 + col) <= 218608) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 218609 && (row * 640 + col) <= 218609) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218610 && (row * 640 + col) <= 218742) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 218743 && (row * 640 + col) <= 218746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218747 && (row * 640 + col) <= 218774) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 218775 && (row * 640 + col) <= 218777) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218778 && (row * 640 + col) <= 218808) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 218809 && (row * 640 + col) <= 218818) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 218819 && (row * 640 + col) <= 219223) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 219224 && (row * 640 + col) <= 219224) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219225 && (row * 640 + col) <= 219248) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 219249 && (row * 640 + col) <= 219249) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219250 && (row * 640 + col) <= 219381) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 219382 && (row * 640 + col) <= 219386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219387 && (row * 640 + col) <= 219414) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 219415 && (row * 640 + col) <= 219417) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219418 && (row * 640 + col) <= 219448) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 219449 && (row * 640 + col) <= 219460) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219461 && (row * 640 + col) <= 219863) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 219864 && (row * 640 + col) <= 219864) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219865 && (row * 640 + col) <= 219888) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 219889 && (row * 640 + col) <= 219889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 219890 && (row * 640 + col) <= 220021) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 220022 && (row * 640 + col) <= 220026) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220027 && (row * 640 + col) <= 220054) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 220055 && (row * 640 + col) <= 220057) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220058 && (row * 640 + col) <= 220088) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 220089 && (row * 640 + col) <= 220100) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220101 && (row * 640 + col) <= 220504) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 220505 && (row * 640 + col) <= 220505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220506 && (row * 640 + col) <= 220527) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 220528 && (row * 640 + col) <= 220528) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220529 && (row * 640 + col) <= 220660) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 220661 && (row * 640 + col) <= 220666) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220667 && (row * 640 + col) <= 220694) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 220695 && (row * 640 + col) <= 220697) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220698 && (row * 640 + col) <= 220728) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 220729 && (row * 640 + col) <= 220745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 220746 && (row * 640 + col) <= 221144) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 221145 && (row * 640 + col) <= 221145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221146 && (row * 640 + col) <= 221149) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 221150 && (row * 640 + col) <= 221161) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221162 && (row * 640 + col) <= 221167) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 221168 && (row * 640 + col) <= 221168) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221169 && (row * 640 + col) <= 221300) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 221301 && (row * 640 + col) <= 221307) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221308 && (row * 640 + col) <= 221334) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 221335 && (row * 640 + col) <= 221337) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221338 && (row * 640 + col) <= 221368) color_data <= 12'b100111011110; else
        if ((row * 640 + col) >= 221369 && (row * 640 + col) <= 221386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221387 && (row * 640 + col) <= 221784) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 221785 && (row * 640 + col) <= 221785) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221786 && (row * 640 + col) <= 221789) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 221790 && (row * 640 + col) <= 221791) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221792 && (row * 640 + col) <= 221799) color_data <= 12'b111011101110; else
        if ((row * 640 + col) >= 221800 && (row * 640 + col) <= 221801) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221802 && (row * 640 + col) <= 221807) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 221808 && (row * 640 + col) <= 221808) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 221809 && (row * 640 + col) <= 221922) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 221923 && (row * 640 + col) <= 222027) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 222028 && (row * 640 + col) <= 222425) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 222426 && (row * 640 + col) <= 222426) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 222427 && (row * 640 + col) <= 222430) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 222431 && (row * 640 + col) <= 222432) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 222433 && (row * 640 + col) <= 222439) color_data <= 12'b111011101110; else
        if ((row * 640 + col) >= 222440 && (row * 640 + col) <= 222440) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 222441 && (row * 640 + col) <= 222446) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 222447 && (row * 640 + col) <= 222447) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 222448 && (row * 640 + col) <= 222559) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 222560 && (row * 640 + col) <= 222668) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 222669 && (row * 640 + col) <= 223066) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 223067 && (row * 640 + col) <= 223067) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223068 && (row * 640 + col) <= 223071) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 223072 && (row * 640 + col) <= 223075) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223076 && (row * 640 + col) <= 223078) color_data <= 12'b111011101110; else
        if ((row * 640 + col) >= 223079 && (row * 640 + col) <= 223080) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223081 && (row * 640 + col) <= 223085) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 223086 && (row * 640 + col) <= 223086) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223087 && (row * 640 + col) <= 223197) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 223198 && (row * 640 + col) <= 223309) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223310 && (row * 640 + col) <= 223706) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 223707 && (row * 640 + col) <= 223707) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223708 && (row * 640 + col) <= 223714) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 223715 && (row * 640 + col) <= 223719) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223720 && (row * 640 + col) <= 223725) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 223726 && (row * 640 + col) <= 223726) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223727 && (row * 640 + col) <= 223834) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 223835 && (row * 640 + col) <= 223951) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 223952 && (row * 640 + col) <= 224347) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 224348 && (row * 640 + col) <= 224349) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 224350 && (row * 640 + col) <= 224363) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 224364 && (row * 640 + col) <= 224365) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 224366 && (row * 640 + col) <= 224469) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 224470 && (row * 640 + col) <= 224507) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 224508 && (row * 640 + col) <= 224534) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 224535 && (row * 640 + col) <= 224537) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 224538 && (row * 640 + col) <= 224567) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 224568 && (row * 640 + col) <= 224593) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 224594 && (row * 640 + col) <= 224989) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 224990 && (row * 640 + col) <= 224990) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 224991 && (row * 640 + col) <= 225002) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 225003 && (row * 640 + col) <= 225003) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 225004 && (row * 640 + col) <= 225107) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 225108 && (row * 640 + col) <= 225122) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 225123 && (row * 640 + col) <= 225144) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225145 && (row * 640 + col) <= 225147) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225148 && (row * 640 + col) <= 225174) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225175 && (row * 640 + col) <= 225177) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225178 && (row * 640 + col) <= 225208) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225209 && (row * 640 + col) <= 225211) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225212 && (row * 640 + col) <= 225221) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225222 && (row * 640 + col) <= 225225) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 225226 && (row * 640 + col) <= 225234) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 225235 && (row * 640 + col) <= 225630) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 225631 && (row * 640 + col) <= 225631) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 225632 && (row * 640 + col) <= 225641) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 225642 && (row * 640 + col) <= 225642) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 225643 && (row * 640 + col) <= 225746) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 225747 && (row * 640 + col) <= 225759) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 225760 && (row * 640 + col) <= 225784) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225785 && (row * 640 + col) <= 225787) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225788 && (row * 640 + col) <= 225803) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225804 && (row * 640 + col) <= 225810) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225811 && (row * 640 + col) <= 225814) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225815 && (row * 640 + col) <= 225817) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225818 && (row * 640 + col) <= 225835) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225836 && (row * 640 + col) <= 225843) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225844 && (row * 640 + col) <= 225848) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225849 && (row * 640 + col) <= 225851) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 225852 && (row * 640 + col) <= 225864) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 225865 && (row * 640 + col) <= 225874) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 225875 && (row * 640 + col) <= 226242) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 226243 && (row * 640 + col) <= 226272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 226273 && (row * 640 + col) <= 226280) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 226281 && (row * 640 + col) <= 226317) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 226318 && (row * 640 + col) <= 226385) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 226386 && (row * 640 + col) <= 226396) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 226397 && (row * 640 + col) <= 226424) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 226425 && (row * 640 + col) <= 226427) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 226428 && (row * 640 + col) <= 226443) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 226444 && (row * 640 + col) <= 226450) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 226451 && (row * 640 + col) <= 226454) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 226455 && (row * 640 + col) <= 226457) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 226458 && (row * 640 + col) <= 226475) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 226476 && (row * 640 + col) <= 226483) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 226484 && (row * 640 + col) <= 226488) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 226489 && (row * 640 + col) <= 226491) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 226492 && (row * 640 + col) <= 226503) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 226504 && (row * 640 + col) <= 226514) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 226515 && (row * 640 + col) <= 226882) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 226883 && (row * 640 + col) <= 226883) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 226884 && (row * 640 + col) <= 226899) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 226900 && (row * 640 + col) <= 226935) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 226936 && (row * 640 + col) <= 226956) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 226957 && (row * 640 + col) <= 226957) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 226958 && (row * 640 + col) <= 227021) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 227022 && (row * 640 + col) <= 227033) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 227034 && (row * 640 + col) <= 227034) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 227035 && (row * 640 + col) <= 227064) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227065 && (row * 640 + col) <= 227067) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227068 && (row * 640 + col) <= 227083) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227084 && (row * 640 + col) <= 227090) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227091 && (row * 640 + col) <= 227094) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227095 && (row * 640 + col) <= 227097) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227098 && (row * 640 + col) <= 227115) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227116 && (row * 640 + col) <= 227123) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227124 && (row * 640 + col) <= 227128) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227129 && (row * 640 + col) <= 227131) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227132 && (row * 640 + col) <= 227143) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227144 && (row * 640 + col) <= 227154) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 227155 && (row * 640 + col) <= 227522) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 227523 && (row * 640 + col) <= 227523) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 227524 && (row * 640 + col) <= 227539) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 227540 && (row * 640 + col) <= 227575) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 227576 && (row * 640 + col) <= 227596) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 227597 && (row * 640 + col) <= 227597) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 227598 && (row * 640 + col) <= 227661) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 227662 && (row * 640 + col) <= 227673) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 227674 && (row * 640 + col) <= 227704) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227705 && (row * 640 + col) <= 227707) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227708 && (row * 640 + col) <= 227734) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227735 && (row * 640 + col) <= 227737) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227738 && (row * 640 + col) <= 227768) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227769 && (row * 640 + col) <= 227771) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 227772 && (row * 640 + col) <= 227782) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 227783 && (row * 640 + col) <= 227796) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 227797 && (row * 640 + col) <= 228162) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 228163 && (row * 640 + col) <= 228163) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 228164 && (row * 640 + col) <= 228179) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 228180 && (row * 640 + col) <= 228215) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 228216 && (row * 640 + col) <= 228236) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 228237 && (row * 640 + col) <= 228237) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 228238 && (row * 640 + col) <= 228300) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 228301 && (row * 640 + col) <= 228313) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 228314 && (row * 640 + col) <= 228344) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 228345 && (row * 640 + col) <= 228347) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 228348 && (row * 640 + col) <= 228374) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 228375 && (row * 640 + col) <= 228377) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 228378 && (row * 640 + col) <= 228408) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 228409 && (row * 640 + col) <= 228411) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 228412 && (row * 640 + col) <= 228422) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 228423 && (row * 640 + col) <= 228436) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 228437 && (row * 640 + col) <= 228802) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 228803 && (row * 640 + col) <= 228803) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 228804 && (row * 640 + col) <= 228819) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 228820 && (row * 640 + col) <= 228855) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 228856 && (row * 640 + col) <= 228876) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 228877 && (row * 640 + col) <= 228877) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 228878 && (row * 640 + col) <= 228940) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 228941 && (row * 640 + col) <= 228953) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 228954 && (row * 640 + col) <= 228984) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 228985 && (row * 640 + col) <= 228987) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 228988 && (row * 640 + col) <= 229014) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 229015 && (row * 640 + col) <= 229017) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 229018 && (row * 640 + col) <= 229048) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 229049 && (row * 640 + col) <= 229051) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 229052 && (row * 640 + col) <= 229062) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 229063 && (row * 640 + col) <= 229076) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 229077 && (row * 640 + col) <= 229442) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 229443 && (row * 640 + col) <= 229443) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 229444 && (row * 640 + col) <= 229459) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 229460 && (row * 640 + col) <= 229495) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 229496 && (row * 640 + col) <= 229516) color_data <= 12'b111111111010; else
        if ((row * 640 + col) >= 229517 && (row * 640 + col) <= 229517) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 229518 && (row * 640 + col) <= 229579) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 229580 && (row * 640 + col) <= 229592) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 229593 && (row * 640 + col) <= 229624) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 229625 && (row * 640 + col) <= 229627) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 229628 && (row * 640 + col) <= 229654) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 229655 && (row * 640 + col) <= 229657) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 229658 && (row * 640 + col) <= 229688) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 229689 && (row * 640 + col) <= 229690) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 229691 && (row * 640 + col) <= 229705) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 229706 && (row * 640 + col) <= 229716) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 229717 && (row * 640 + col) <= 230082) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 230083 && (row * 640 + col) <= 230105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 230106 && (row * 640 + col) <= 230129) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 230130 && (row * 640 + col) <= 230157) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 230158 && (row * 640 + col) <= 230219) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 230220 && (row * 640 + col) <= 230231) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 230232 && (row * 640 + col) <= 230264) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230265 && (row * 640 + col) <= 230267) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 230268 && (row * 640 + col) <= 230294) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230295 && (row * 640 + col) <= 230297) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 230298 && (row * 640 + col) <= 230327) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230328 && (row * 640 + col) <= 230330) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 230331 && (row * 640 + col) <= 230345) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230346 && (row * 640 + col) <= 230356) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 230357 && (row * 640 + col) <= 230744) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 230745 && (row * 640 + col) <= 230745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 230746 && (row * 640 + col) <= 230769) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 230770 && (row * 640 + col) <= 230770) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 230771 && (row * 640 + col) <= 230859) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 230860 && (row * 640 + col) <= 230871) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 230872 && (row * 640 + col) <= 230904) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230905 && (row * 640 + col) <= 230907) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 230908 && (row * 640 + col) <= 230934) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230935 && (row * 640 + col) <= 230937) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 230938 && (row * 640 + col) <= 230967) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230968 && (row * 640 + col) <= 230970) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 230971 && (row * 640 + col) <= 230985) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 230986 && (row * 640 + col) <= 230996) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 230997 && (row * 640 + col) <= 231384) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 231385 && (row * 640 + col) <= 231385) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 231386 && (row * 640 + col) <= 231409) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 231410 && (row * 640 + col) <= 231410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 231411 && (row * 640 + col) <= 231499) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 231500 && (row * 640 + col) <= 231509) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 231510 && (row * 640 + col) <= 231544) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 231545 && (row * 640 + col) <= 231547) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 231548 && (row * 640 + col) <= 231574) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 231575 && (row * 640 + col) <= 231577) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 231578 && (row * 640 + col) <= 231607) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 231608 && (row * 640 + col) <= 231610) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 231611 && (row * 640 + col) <= 231627) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 231628 && (row * 640 + col) <= 231632) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 231633 && (row * 640 + col) <= 231636) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 231637 && (row * 640 + col) <= 232024) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 232025 && (row * 640 + col) <= 232025) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 232026 && (row * 640 + col) <= 232049) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 232050 && (row * 640 + col) <= 232050) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 232051 && (row * 640 + col) <= 232139) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 232140 && (row * 640 + col) <= 232148) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 232149 && (row * 640 + col) <= 232184) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232185 && (row * 640 + col) <= 232187) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 232188 && (row * 640 + col) <= 232214) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232215 && (row * 640 + col) <= 232217) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 232218 && (row * 640 + col) <= 232247) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232248 && (row * 640 + col) <= 232250) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 232251 && (row * 640 + col) <= 232267) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232268 && (row * 640 + col) <= 232274) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 232275 && (row * 640 + col) <= 232664) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 232665 && (row * 640 + col) <= 232665) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 232666 && (row * 640 + col) <= 232689) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 232690 && (row * 640 + col) <= 232690) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 232691 && (row * 640 + col) <= 232779) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 232780 && (row * 640 + col) <= 232787) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 232788 && (row * 640 + col) <= 232824) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232825 && (row * 640 + col) <= 232827) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 232828 && (row * 640 + col) <= 232854) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232855 && (row * 640 + col) <= 232857) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 232858 && (row * 640 + col) <= 232885) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232886 && (row * 640 + col) <= 232890) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 232891 && (row * 640 + col) <= 232907) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 232908 && (row * 640 + col) <= 232914) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 232915 && (row * 640 + col) <= 233304) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 233305 && (row * 640 + col) <= 233305) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 233306 && (row * 640 + col) <= 233329) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 233330 && (row * 640 + col) <= 233330) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 233331 && (row * 640 + col) <= 233418) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 233419 && (row * 640 + col) <= 233422) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 233423 && (row * 640 + col) <= 233425) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 233426 && (row * 640 + col) <= 233464) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 233465 && (row * 640 + col) <= 233467) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 233468 && (row * 640 + col) <= 233494) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 233495 && (row * 640 + col) <= 233497) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 233498 && (row * 640 + col) <= 233522) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 233523 && (row * 640 + col) <= 233530) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 233531 && (row * 640 + col) <= 233547) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 233548 && (row * 640 + col) <= 233554) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 233555 && (row * 640 + col) <= 233944) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 233945 && (row * 640 + col) <= 233945) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 233946 && (row * 640 + col) <= 233969) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 233970 && (row * 640 + col) <= 233970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 233971 && (row * 640 + col) <= 234058) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 234059 && (row * 640 + col) <= 234065) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 234066 && (row * 640 + col) <= 234104) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234105 && (row * 640 + col) <= 234107) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 234108 && (row * 640 + col) <= 234134) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234135 && (row * 640 + col) <= 234137) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 234138 && (row * 640 + col) <= 234160) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234161 && (row * 640 + col) <= 234170) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 234171 && (row * 640 + col) <= 234187) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234188 && (row * 640 + col) <= 234194) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 234195 && (row * 640 + col) <= 234584) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 234585 && (row * 640 + col) <= 234585) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 234586 && (row * 640 + col) <= 234609) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 234610 && (row * 640 + col) <= 234610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 234611 && (row * 640 + col) <= 234697) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 234698 && (row * 640 + col) <= 234704) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 234705 && (row * 640 + col) <= 234744) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234745 && (row * 640 + col) <= 234747) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 234748 && (row * 640 + col) <= 234774) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234775 && (row * 640 + col) <= 234777) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 234778 && (row * 640 + col) <= 234797) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234798 && (row * 640 + col) <= 234805) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 234806 && (row * 640 + col) <= 234827) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 234828 && (row * 640 + col) <= 234834) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 234835 && (row * 640 + col) <= 235224) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 235225 && (row * 640 + col) <= 235225) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 235226 && (row * 640 + col) <= 235249) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 235250 && (row * 640 + col) <= 235250) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 235251 && (row * 640 + col) <= 235337) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 235338 && (row * 640 + col) <= 235344) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 235345 && (row * 640 + col) <= 235384) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 235385 && (row * 640 + col) <= 235387) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 235388 && (row * 640 + col) <= 235414) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 235415 && (row * 640 + col) <= 235417) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 235418 && (row * 640 + col) <= 235435) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 235436 && (row * 640 + col) <= 235443) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 235444 && (row * 640 + col) <= 235467) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 235468 && (row * 640 + col) <= 235474) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 235475 && (row * 640 + col) <= 235864) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 235865 && (row * 640 + col) <= 235865) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 235866 && (row * 640 + col) <= 235889) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 235890 && (row * 640 + col) <= 235890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 235891 && (row * 640 + col) <= 235977) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 235978 && (row * 640 + col) <= 235983) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 235984 && (row * 640 + col) <= 236024) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236025 && (row * 640 + col) <= 236027) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 236028 && (row * 640 + col) <= 236054) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236055 && (row * 640 + col) <= 236057) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 236058 && (row * 640 + col) <= 236072) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236073 && (row * 640 + col) <= 236080) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 236081 && (row * 640 + col) <= 236107) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236108 && (row * 640 + col) <= 236114) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 236115 && (row * 640 + col) <= 236504) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 236505 && (row * 640 + col) <= 236505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 236506 && (row * 640 + col) <= 236529) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 236530 && (row * 640 + col) <= 236530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 236531 && (row * 640 + col) <= 236617) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 236618 && (row * 640 + col) <= 236623) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 236624 && (row * 640 + col) <= 236649) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236650 && (row * 640 + col) <= 236656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 236657 && (row * 640 + col) <= 236664) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236665 && (row * 640 + col) <= 236667) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 236668 && (row * 640 + col) <= 236694) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236695 && (row * 640 + col) <= 236697) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 236698 && (row * 640 + col) <= 236710) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236711 && (row * 640 + col) <= 236718) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 236719 && (row * 640 + col) <= 236724) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 236725 && (row * 640 + col) <= 236747) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 236748 && (row * 640 + col) <= 236754) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 236755 && (row * 640 + col) <= 237144) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 237145 && (row * 640 + col) <= 237145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237146 && (row * 640 + col) <= 237169) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 237170 && (row * 640 + col) <= 237170) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237171 && (row * 640 + col) <= 237257) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 237258 && (row * 640 + col) <= 237263) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237264 && (row * 640 + col) <= 237287) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 237288 && (row * 640 + col) <= 237298) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237299 && (row * 640 + col) <= 237304) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 237305 && (row * 640 + col) <= 237307) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 237308 && (row * 640 + col) <= 237334) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 237335 && (row * 640 + col) <= 237337) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 237338 && (row * 640 + col) <= 237347) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 237348 && (row * 640 + col) <= 237356) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 237357 && (row * 640 + col) <= 237366) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237367 && (row * 640 + col) <= 237387) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 237388 && (row * 640 + col) <= 237393) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237394 && (row * 640 + col) <= 237784) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 237785 && (row * 640 + col) <= 237785) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237786 && (row * 640 + col) <= 237809) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 237810 && (row * 640 + col) <= 237810) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237811 && (row * 640 + col) <= 237897) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 237898 && (row * 640 + col) <= 237903) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237904 && (row * 640 + col) <= 237925) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 237926 && (row * 640 + col) <= 237940) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 237941 && (row * 640 + col) <= 237993) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 237994 && (row * 640 + col) <= 238008) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238009 && (row * 640 + col) <= 238027) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 238028 && (row * 640 + col) <= 238033) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238034 && (row * 640 + col) <= 238424) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 238425 && (row * 640 + col) <= 238425) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238426 && (row * 640 + col) <= 238449) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 238450 && (row * 640 + col) <= 238450) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238451 && (row * 640 + col) <= 238537) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 238538 && (row * 640 + col) <= 238543) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238544 && (row * 640 + col) <= 238565) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 238566 && (row * 640 + col) <= 238580) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238581 && (row * 640 + col) <= 238632) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 238633 && (row * 640 + col) <= 238648) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238649 && (row * 640 + col) <= 238667) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 238668 && (row * 640 + col) <= 238673) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 238674 && (row * 640 + col) <= 239064) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 239065 && (row * 640 + col) <= 239065) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239066 && (row * 640 + col) <= 239089) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 239090 && (row * 640 + col) <= 239090) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239091 && (row * 640 + col) <= 239177) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 239178 && (row * 640 + col) <= 239183) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239184 && (row * 640 + col) <= 239205) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 239206 && (row * 640 + col) <= 239220) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239221 && (row * 640 + col) <= 239272) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 239273 && (row * 640 + col) <= 239288) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239289 && (row * 640 + col) <= 239307) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 239308 && (row * 640 + col) <= 239312) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239313 && (row * 640 + col) <= 239704) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 239705 && (row * 640 + col) <= 239705) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239706 && (row * 640 + col) <= 239729) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 239730 && (row * 640 + col) <= 239730) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239731 && (row * 640 + col) <= 239817) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 239818 && (row * 640 + col) <= 239824) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239825 && (row * 640 + col) <= 239842) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 239843 && (row * 640 + col) <= 239863) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239864 && (row * 640 + col) <= 239864) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 239865 && (row * 640 + col) <= 239867) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 239868 && (row * 640 + col) <= 239894) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 239895 && (row * 640 + col) <= 239897) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 239898 && (row * 640 + col) <= 239907) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 239908 && (row * 640 + col) <= 239910) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 239911 && (row * 640 + col) <= 239931) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239932 && (row * 640 + col) <= 239946) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 239947 && (row * 640 + col) <= 239952) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 239953 && (row * 640 + col) <= 239999) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240000 && (row * 640 + col) <= 240049) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240050 && (row * 640 + col) <= 240100) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240101 && (row * 640 + col) <= 240149) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240150 && (row * 640 + col) <= 240200) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240201 && (row * 640 + col) <= 240249) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240250 && (row * 640 + col) <= 240300) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240301 && (row * 640 + col) <= 240344) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240345 && (row * 640 + col) <= 240345) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240346 && (row * 640 + col) <= 240369) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 240370 && (row * 640 + col) <= 240370) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240371 && (row * 640 + col) <= 240400) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240401 && (row * 640 + col) <= 240449) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240450 && (row * 640 + col) <= 240458) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240459 && (row * 640 + col) <= 240465) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240466 && (row * 640 + col) <= 240482) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 240483 && (row * 640 + col) <= 240503) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240504 && (row * 640 + col) <= 240504) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 240505 && (row * 640 + col) <= 240507) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 240508 && (row * 640 + col) <= 240534) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 240535 && (row * 640 + col) <= 240537) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 240538 && (row * 640 + col) <= 240547) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 240548 && (row * 640 + col) <= 240550) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 240551 && (row * 640 + col) <= 240571) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240572 && (row * 640 + col) <= 240586) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 240587 && (row * 640 + col) <= 240592) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240593 && (row * 640 + col) <= 240600) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240601 && (row * 640 + col) <= 240689) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240690 && (row * 640 + col) <= 240740) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240741 && (row * 640 + col) <= 240789) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240790 && (row * 640 + col) <= 240840) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240841 && (row * 640 + col) <= 240889) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240890 && (row * 640 + col) <= 240940) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 240941 && (row * 640 + col) <= 240984) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 240985 && (row * 640 + col) <= 240985) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 240986 && (row * 640 + col) <= 241009) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 241010 && (row * 640 + col) <= 241010) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241011 && (row * 640 + col) <= 241040) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241041 && (row * 640 + col) <= 241089) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241090 && (row * 640 + col) <= 241098) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241099 && (row * 640 + col) <= 241105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241106 && (row * 640 + col) <= 241121) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 241122 && (row * 640 + col) <= 241130) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241131 && (row * 640 + col) <= 241135) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 241136 && (row * 640 + col) <= 241144) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241145 && (row * 640 + col) <= 241149) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 241150 && (row * 640 + col) <= 241174) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 241175 && (row * 640 + col) <= 241177) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 241178 && (row * 640 + col) <= 241187) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 241188 && (row * 640 + col) <= 241190) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 241191 && (row * 640 + col) <= 241198) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241199 && (row * 640 + col) <= 241203) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 241204 && (row * 640 + col) <= 241212) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241213 && (row * 640 + col) <= 241226) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 241227 && (row * 640 + col) <= 241232) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241233 && (row * 640 + col) <= 241240) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241241 && (row * 640 + col) <= 241329) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241330 && (row * 640 + col) <= 241380) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241381 && (row * 640 + col) <= 241429) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241430 && (row * 640 + col) <= 241480) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241481 && (row * 640 + col) <= 241529) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241530 && (row * 640 + col) <= 241580) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241581 && (row * 640 + col) <= 241624) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241625 && (row * 640 + col) <= 241625) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241626 && (row * 640 + col) <= 241649) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 241650 && (row * 640 + col) <= 241650) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241651 && (row * 640 + col) <= 241680) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241681 && (row * 640 + col) <= 241729) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241730 && (row * 640 + col) <= 241738) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241739 && (row * 640 + col) <= 241747) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241748 && (row * 640 + col) <= 241761) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 241762 && (row * 640 + col) <= 241769) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241770 && (row * 640 + col) <= 241776) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 241777 && (row * 640 + col) <= 241784) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241785 && (row * 640 + col) <= 241830) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 241831 && (row * 640 + col) <= 241837) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241838 && (row * 640 + col) <= 241844) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 241845 && (row * 640 + col) <= 241852) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241853 && (row * 640 + col) <= 241865) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 241866 && (row * 640 + col) <= 241871) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 241872 && (row * 640 + col) <= 241880) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 241881 && (row * 640 + col) <= 241969) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 241970 && (row * 640 + col) <= 242020) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242021 && (row * 640 + col) <= 242069) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242070 && (row * 640 + col) <= 242120) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242121 && (row * 640 + col) <= 242169) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242170 && (row * 640 + col) <= 242220) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242221 && (row * 640 + col) <= 242264) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242265 && (row * 640 + col) <= 242265) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242266 && (row * 640 + col) <= 242289) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 242290 && (row * 640 + col) <= 242290) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242291 && (row * 640 + col) <= 242320) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242321 && (row * 640 + col) <= 242369) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242370 && (row * 640 + col) <= 242379) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242380 && (row * 640 + col) <= 242389) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242390 && (row * 640 + col) <= 242400) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 242401 && (row * 640 + col) <= 242408) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242409 && (row * 640 + col) <= 242417) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 242418 && (row * 640 + col) <= 242425) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242426 && (row * 640 + col) <= 242426) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 242427 && (row * 640 + col) <= 242468) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 242469 && (row * 640 + col) <= 242476) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242477 && (row * 640 + col) <= 242485) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 242486 && (row * 640 + col) <= 242493) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242494 && (row * 640 + col) <= 242505) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 242506 && (row * 640 + col) <= 242511) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242512 && (row * 640 + col) <= 242520) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242521 && (row * 640 + col) <= 242609) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242610 && (row * 640 + col) <= 242660) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242661 && (row * 640 + col) <= 242709) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242710 && (row * 640 + col) <= 242760) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242761 && (row * 640 + col) <= 242809) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242810 && (row * 640 + col) <= 242860) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242861 && (row * 640 + col) <= 242904) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 242905 && (row * 640 + col) <= 242905) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242906 && (row * 640 + col) <= 242929) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 242930 && (row * 640 + col) <= 242930) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 242931 && (row * 640 + col) <= 242960) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 242961 && (row * 640 + col) <= 243009) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243010 && (row * 640 + col) <= 243019) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243020 && (row * 640 + col) <= 243030) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243031 && (row * 640 + col) <= 243040) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 243041 && (row * 640 + col) <= 243047) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243048 && (row * 640 + col) <= 243058) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 243059 && (row * 640 + col) <= 243065) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243066 && (row * 640 + col) <= 243066) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 243067 && (row * 640 + col) <= 243108) color_data <= 12'b001101110010; else
        if ((row * 640 + col) >= 243109 && (row * 640 + col) <= 243115) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243116 && (row * 640 + col) <= 243126) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 243127 && (row * 640 + col) <= 243133) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243134 && (row * 640 + col) <= 243144) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 243145 && (row * 640 + col) <= 243150) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243151 && (row * 640 + col) <= 243160) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243161 && (row * 640 + col) <= 243249) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243250 && (row * 640 + col) <= 243300) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243301 && (row * 640 + col) <= 243349) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243350 && (row * 640 + col) <= 243400) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243401 && (row * 640 + col) <= 243449) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243450 && (row * 640 + col) <= 243500) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243501 && (row * 640 + col) <= 243544) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243545 && (row * 640 + col) <= 243545) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243546 && (row * 640 + col) <= 243569) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 243570 && (row * 640 + col) <= 243570) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243571 && (row * 640 + col) <= 243600) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243601 && (row * 640 + col) <= 243649) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243650 && (row * 640 + col) <= 243660) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243661 && (row * 640 + col) <= 243673) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243674 && (row * 640 + col) <= 243680) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 243681 && (row * 640 + col) <= 243687) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243688 && (row * 640 + col) <= 243698) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 243699 && (row * 640 + col) <= 243705) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243706 && (row * 640 + col) <= 243748) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 243749 && (row * 640 + col) <= 243755) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243756 && (row * 640 + col) <= 243766) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 243767 && (row * 640 + col) <= 243773) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243774 && (row * 640 + col) <= 243783) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 243784 && (row * 640 + col) <= 243789) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 243790 && (row * 640 + col) <= 243800) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243801 && (row * 640 + col) <= 243889) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243890 && (row * 640 + col) <= 243940) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 243941 && (row * 640 + col) <= 243989) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 243990 && (row * 640 + col) <= 244040) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244041 && (row * 640 + col) <= 244089) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244090 && (row * 640 + col) <= 244140) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244141 && (row * 640 + col) <= 244184) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244185 && (row * 640 + col) <= 244185) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244186 && (row * 640 + col) <= 244209) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 244210 && (row * 640 + col) <= 244210) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244211 && (row * 640 + col) <= 244240) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244241 && (row * 640 + col) <= 244289) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244290 && (row * 640 + col) <= 244303) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244304 && (row * 640 + col) <= 244316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244317 && (row * 640 + col) <= 244320) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 244321 && (row * 640 + col) <= 244327) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244328 && (row * 640 + col) <= 244338) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 244339 && (row * 640 + col) <= 244345) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244346 && (row * 640 + col) <= 244388) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 244389 && (row * 640 + col) <= 244395) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244396 && (row * 640 + col) <= 244406) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 244407 && (row * 640 + col) <= 244413) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244414 && (row * 640 + col) <= 244419) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 244420 && (row * 640 + col) <= 244428) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244429 && (row * 640 + col) <= 244440) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244441 && (row * 640 + col) <= 244529) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244530 && (row * 640 + col) <= 244580) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244581 && (row * 640 + col) <= 244629) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244630 && (row * 640 + col) <= 244680) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244681 && (row * 640 + col) <= 244729) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244730 && (row * 640 + col) <= 244780) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244781 && (row * 640 + col) <= 244824) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244825 && (row * 640 + col) <= 244825) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244826 && (row * 640 + col) <= 244849) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 244850 && (row * 640 + col) <= 244850) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244851 && (row * 640 + col) <= 244880) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244881 && (row * 640 + col) <= 244929) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 244930 && (row * 640 + col) <= 244944) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 244945 && (row * 640 + col) <= 244967) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 244968 && (row * 640 + col) <= 244978) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 244979 && (row * 640 + col) <= 245035) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245036 && (row * 640 + col) <= 245046) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 245047 && (row * 640 + col) <= 245067) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245068 && (row * 640 + col) <= 245080) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245081 && (row * 640 + col) <= 245169) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245170 && (row * 640 + col) <= 245220) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245221 && (row * 640 + col) <= 245269) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245270 && (row * 640 + col) <= 245320) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245321 && (row * 640 + col) <= 245369) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245370 && (row * 640 + col) <= 245420) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245421 && (row * 640 + col) <= 245464) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245465 && (row * 640 + col) <= 245465) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245466 && (row * 640 + col) <= 245489) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 245490 && (row * 640 + col) <= 245490) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245491 && (row * 640 + col) <= 245520) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245521 && (row * 640 + col) <= 245569) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245570 && (row * 640 + col) <= 245585) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245586 && (row * 640 + col) <= 245607) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245608 && (row * 640 + col) <= 245618) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 245619 && (row * 640 + col) <= 245675) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245676 && (row * 640 + col) <= 245686) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 245687 && (row * 640 + col) <= 245706) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 245707 && (row * 640 + col) <= 245720) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245721 && (row * 640 + col) <= 245809) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245810 && (row * 640 + col) <= 245860) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245861 && (row * 640 + col) <= 245909) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 245910 && (row * 640 + col) <= 245960) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 245961 && (row * 640 + col) <= 246009) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246010 && (row * 640 + col) <= 246060) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246061 && (row * 640 + col) <= 246104) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246105 && (row * 640 + col) <= 246105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246106 && (row * 640 + col) <= 246129) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 246130 && (row * 640 + col) <= 246130) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246131 && (row * 640 + col) <= 246160) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246161 && (row * 640 + col) <= 246209) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246210 && (row * 640 + col) <= 246227) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246228 && (row * 640 + col) <= 246248) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246249 && (row * 640 + col) <= 246257) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 246258 && (row * 640 + col) <= 246316) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246317 && (row * 640 + col) <= 246325) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 246326 && (row * 640 + col) <= 246345) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246346 && (row * 640 + col) <= 246360) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246361 && (row * 640 + col) <= 246449) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246450 && (row * 640 + col) <= 246500) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246501 && (row * 640 + col) <= 246549) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246550 && (row * 640 + col) <= 246600) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246601 && (row * 640 + col) <= 246649) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246650 && (row * 640 + col) <= 246700) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246701 && (row * 640 + col) <= 246744) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246745 && (row * 640 + col) <= 246745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246746 && (row * 640 + col) <= 246769) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 246770 && (row * 640 + col) <= 246770) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246771 && (row * 640 + col) <= 246800) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246801 && (row * 640 + col) <= 246849) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 246850 && (row * 640 + col) <= 246868) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 246869 && (row * 640 + col) <= 246889) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246890 && (row * 640 + col) <= 246896) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 246897 && (row * 640 + col) <= 246957) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246958 && (row * 640 + col) <= 246964) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 246965 && (row * 640 + col) <= 246984) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 246985 && (row * 640 + col) <= 247000) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247001 && (row * 640 + col) <= 247089) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247090 && (row * 640 + col) <= 247140) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247141 && (row * 640 + col) <= 247189) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247190 && (row * 640 + col) <= 247240) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247241 && (row * 640 + col) <= 247289) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247290 && (row * 640 + col) <= 247340) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247341 && (row * 640 + col) <= 247384) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247385 && (row * 640 + col) <= 247385) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247386 && (row * 640 + col) <= 247409) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 247410 && (row * 640 + col) <= 247410) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247411 && (row * 640 + col) <= 247440) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247441 && (row * 640 + col) <= 247489) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247490 && (row * 640 + col) <= 247512) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247513 && (row * 640 + col) <= 247530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247531 && (row * 640 + col) <= 247535) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 247536 && (row * 640 + col) <= 247598) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247599 && (row * 640 + col) <= 247603) color_data <= 12'b011101110111; else
        if ((row * 640 + col) >= 247604 && (row * 640 + col) <= 247621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 247622 && (row * 640 + col) <= 247640) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247641 && (row * 640 + col) <= 247729) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247730 && (row * 640 + col) <= 247780) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247781 && (row * 640 + col) <= 247829) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247830 && (row * 640 + col) <= 247880) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247881 && (row * 640 + col) <= 247929) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 247930 && (row * 640 + col) <= 247980) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 247981 && (row * 640 + col) <= 248024) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248025 && (row * 640 + col) <= 248025) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248026 && (row * 640 + col) <= 248049) color_data <= 12'b111000010010; else
        if ((row * 640 + col) >= 248050 && (row * 640 + col) <= 248050) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248051 && (row * 640 + col) <= 248080) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248081 && (row * 640 + col) <= 248129) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248130 && (row * 640 + col) <= 248155) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248156 && (row * 640 + col) <= 248183) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248184 && (row * 640 + col) <= 248230) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248231 && (row * 640 + col) <= 248257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248258 && (row * 640 + col) <= 248280) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248281 && (row * 640 + col) <= 248369) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248370 && (row * 640 + col) <= 248420) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248421 && (row * 640 + col) <= 248469) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248470 && (row * 640 + col) <= 248520) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248521 && (row * 640 + col) <= 248569) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248570 && (row * 640 + col) <= 248620) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248621 && (row * 640 + col) <= 248664) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248665 && (row * 640 + col) <= 248665) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248666 && (row * 640 + col) <= 248689) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 248690 && (row * 640 + col) <= 248690) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248691 && (row * 640 + col) <= 248720) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248721 && (row * 640 + col) <= 248769) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248770 && (row * 640 + col) <= 248802) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248803 && (row * 640 + col) <= 248823) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248824 && (row * 640 + col) <= 248870) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248871 && (row * 640 + col) <= 248891) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 248892 && (row * 640 + col) <= 248920) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 248921 && (row * 640 + col) <= 248959) color_data <= 12'b110011001100; else
        if ((row * 640 + col) >= 248960 && (row * 640 + col) <= 249304) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249305 && (row * 640 + col) <= 249305) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249306 && (row * 640 + col) <= 249329) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 249330 && (row * 640 + col) <= 249330) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249331 && (row * 640 + col) <= 249443) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249444 && (row * 640 + col) <= 249462) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249463 && (row * 640 + col) <= 249511) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249512 && (row * 640 + col) <= 249530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249531 && (row * 640 + col) <= 249944) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 249945 && (row * 640 + col) <= 249945) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249946 && (row * 640 + col) <= 249969) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 249970 && (row * 640 + col) <= 249970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249971 && (row * 640 + col) <= 250084) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 250085 && (row * 640 + col) <= 250101) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250102 && (row * 640 + col) <= 250152) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 250153 && (row * 640 + col) <= 250169) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250170 && (row * 640 + col) <= 250584) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 250585 && (row * 640 + col) <= 250585) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250586 && (row * 640 + col) <= 250609) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 250610 && (row * 640 + col) <= 250610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250611 && (row * 640 + col) <= 250725) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 250726 && (row * 640 + col) <= 250740) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250741 && (row * 640 + col) <= 250793) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 250794 && (row * 640 + col) <= 250808) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250809 && (row * 640 + col) <= 251224) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251225 && (row * 640 + col) <= 251225) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251226 && (row * 640 + col) <= 251249) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 251250 && (row * 640 + col) <= 251250) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251251 && (row * 640 + col) <= 251367) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251368 && (row * 640 + col) <= 251378) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251379 && (row * 640 + col) <= 251435) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251436 && (row * 640 + col) <= 251446) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251447 && (row * 640 + col) <= 251864) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 251865 && (row * 640 + col) <= 251865) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251866 && (row * 640 + col) <= 251871) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 251872 && (row * 640 + col) <= 251883) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251884 && (row * 640 + col) <= 251889) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 251890 && (row * 640 + col) <= 251890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251891 && (row * 640 + col) <= 252009) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 252010 && (row * 640 + col) <= 252016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252017 && (row * 640 + col) <= 252077) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 252078 && (row * 640 + col) <= 252084) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252085 && (row * 640 + col) <= 252504) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 252505 && (row * 640 + col) <= 252505) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252506 && (row * 640 + col) <= 252511) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 252512 && (row * 640 + col) <= 252512) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252513 && (row * 640 + col) <= 252522) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 252523 && (row * 640 + col) <= 252523) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252524 && (row * 640 + col) <= 252529) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 252530 && (row * 640 + col) <= 252530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252531 && (row * 640 + col) <= 253144) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 253145 && (row * 640 + col) <= 253145) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253146 && (row * 640 + col) <= 253151) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 253152 && (row * 640 + col) <= 253152) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253153 && (row * 640 + col) <= 253162) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 253163 && (row * 640 + col) <= 253163) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253164 && (row * 640 + col) <= 253169) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 253170 && (row * 640 + col) <= 253170) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253171 && (row * 640 + col) <= 253784) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 253785 && (row * 640 + col) <= 253785) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253786 && (row * 640 + col) <= 253791) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 253792 && (row * 640 + col) <= 253792) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253793 && (row * 640 + col) <= 253802) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 253803 && (row * 640 + col) <= 253803) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253804 && (row * 640 + col) <= 253809) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 253810 && (row * 640 + col) <= 253810) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253811 && (row * 640 + col) <= 254424) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 254425 && (row * 640 + col) <= 254425) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254426 && (row * 640 + col) <= 254431) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 254432 && (row * 640 + col) <= 254432) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254433 && (row * 640 + col) <= 254442) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 254443 && (row * 640 + col) <= 254443) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254444 && (row * 640 + col) <= 254449) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 254450 && (row * 640 + col) <= 254450) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254451 && (row * 640 + col) <= 255064) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 255065 && (row * 640 + col) <= 255065) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255066 && (row * 640 + col) <= 255071) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 255072 && (row * 640 + col) <= 255072) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255073 && (row * 640 + col) <= 255082) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 255083 && (row * 640 + col) <= 255083) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255084 && (row * 640 + col) <= 255089) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 255090 && (row * 640 + col) <= 255090) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255091 && (row * 640 + col) <= 255704) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 255705 && (row * 640 + col) <= 255705) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255706 && (row * 640 + col) <= 255711) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 255712 && (row * 640 + col) <= 255712) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255713 && (row * 640 + col) <= 255722) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 255723 && (row * 640 + col) <= 255723) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255724 && (row * 640 + col) <= 255729) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 255730 && (row * 640 + col) <= 255730) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255731 && (row * 640 + col) <= 256344) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 256345 && (row * 640 + col) <= 256345) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256346 && (row * 640 + col) <= 256351) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 256352 && (row * 640 + col) <= 256352) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256353 && (row * 640 + col) <= 256362) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 256363 && (row * 640 + col) <= 256363) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256364 && (row * 640 + col) <= 256369) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 256370 && (row * 640 + col) <= 256370) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256371 && (row * 640 + col) <= 256984) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 256985 && (row * 640 + col) <= 256985) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256986 && (row * 640 + col) <= 256991) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 256992 && (row * 640 + col) <= 256992) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256993 && (row * 640 + col) <= 257002) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 257003 && (row * 640 + col) <= 257003) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257004 && (row * 640 + col) <= 257009) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 257010 && (row * 640 + col) <= 257010) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257011 && (row * 640 + col) <= 257624) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 257625 && (row * 640 + col) <= 257625) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257626 && (row * 640 + col) <= 257631) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 257632 && (row * 640 + col) <= 257632) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257633 && (row * 640 + col) <= 257642) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 257643 && (row * 640 + col) <= 257643) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257644 && (row * 640 + col) <= 257649) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 257650 && (row * 640 + col) <= 257650) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257651 && (row * 640 + col) <= 258264) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 258265 && (row * 640 + col) <= 258265) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258266 && (row * 640 + col) <= 258271) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 258272 && (row * 640 + col) <= 258272) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258273 && (row * 640 + col) <= 258282) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 258283 && (row * 640 + col) <= 258283) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258284 && (row * 640 + col) <= 258289) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 258290 && (row * 640 + col) <= 258290) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258291 && (row * 640 + col) <= 258904) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 258905 && (row * 640 + col) <= 258905) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258906 && (row * 640 + col) <= 258911) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 258912 && (row * 640 + col) <= 258912) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258913 && (row * 640 + col) <= 258922) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 258923 && (row * 640 + col) <= 258923) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258924 && (row * 640 + col) <= 258929) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 258930 && (row * 640 + col) <= 258930) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 258931 && (row * 640 + col) <= 259544) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 259545 && (row * 640 + col) <= 259545) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259546 && (row * 640 + col) <= 259551) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 259552 && (row * 640 + col) <= 259552) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259553 && (row * 640 + col) <= 259562) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 259563 && (row * 640 + col) <= 259563) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259564 && (row * 640 + col) <= 259569) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 259570 && (row * 640 + col) <= 259570) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 259571 && (row * 640 + col) <= 260184) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 260185 && (row * 640 + col) <= 260185) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260186 && (row * 640 + col) <= 260191) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 260192 && (row * 640 + col) <= 260192) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260193 && (row * 640 + col) <= 260202) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 260203 && (row * 640 + col) <= 260203) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260204 && (row * 640 + col) <= 260209) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 260210 && (row * 640 + col) <= 260210) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260211 && (row * 640 + col) <= 260824) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 260825 && (row * 640 + col) <= 260825) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260826 && (row * 640 + col) <= 260831) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 260832 && (row * 640 + col) <= 260832) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260833 && (row * 640 + col) <= 260842) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 260843 && (row * 640 + col) <= 260843) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260844 && (row * 640 + col) <= 260849) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 260850 && (row * 640 + col) <= 260850) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 260851 && (row * 640 + col) <= 261464) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 261465 && (row * 640 + col) <= 261465) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261466 && (row * 640 + col) <= 261471) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 261472 && (row * 640 + col) <= 261472) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261473 && (row * 640 + col) <= 261482) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 261483 && (row * 640 + col) <= 261483) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261484 && (row * 640 + col) <= 261489) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 261490 && (row * 640 + col) <= 261490) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 261491 && (row * 640 + col) <= 262104) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 262105 && (row * 640 + col) <= 262105) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262106 && (row * 640 + col) <= 262111) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 262112 && (row * 640 + col) <= 262112) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262113 && (row * 640 + col) <= 262122) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 262123 && (row * 640 + col) <= 262123) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262124 && (row * 640 + col) <= 262129) color_data <= 12'b001101001100; else
        if ((row * 640 + col) >= 262130 && (row * 640 + col) <= 262130) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262131 && (row * 640 + col) <= 262735) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 262736 && (row * 640 + col) <= 262745) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262746 && (row * 640 + col) <= 262751) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 262752 && (row * 640 + col) <= 262752) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262753 && (row * 640 + col) <= 262762) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 262763 && (row * 640 + col) <= 262763) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262764 && (row * 640 + col) <= 262769) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 262770 && (row * 640 + col) <= 262781) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 262782 && (row * 640 + col) <= 263375) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 263376 && (row * 640 + col) <= 263376) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263377 && (row * 640 + col) <= 263391) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 263392 && (row * 640 + col) <= 263392) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263393 && (row * 640 + col) <= 263402) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 263403 && (row * 640 + col) <= 263403) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263404 && (row * 640 + col) <= 263420) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 263421 && (row * 640 + col) <= 263421) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 263422 && (row * 640 + col) <= 264015) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 264016 && (row * 640 + col) <= 264016) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264017 && (row * 640 + col) <= 264031) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 264032 && (row * 640 + col) <= 264032) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264033 && (row * 640 + col) <= 264042) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 264043 && (row * 640 + col) <= 264043) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264044 && (row * 640 + col) <= 264060) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 264061 && (row * 640 + col) <= 264061) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264062 && (row * 640 + col) <= 264655) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 264656 && (row * 640 + col) <= 264656) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264657 && (row * 640 + col) <= 264671) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 264672 && (row * 640 + col) <= 264672) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264673 && (row * 640 + col) <= 264682) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 264683 && (row * 640 + col) <= 264683) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264684 && (row * 640 + col) <= 264700) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 264701 && (row * 640 + col) <= 264701) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 264702 && (row * 640 + col) <= 265295) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 265296 && (row * 640 + col) <= 265296) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265297 && (row * 640 + col) <= 265311) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 265312 && (row * 640 + col) <= 265312) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265313 && (row * 640 + col) <= 265322) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 265323 && (row * 640 + col) <= 265323) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265324 && (row * 640 + col) <= 265340) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 265341 && (row * 640 + col) <= 265341) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265342 && (row * 640 + col) <= 265935) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 265936 && (row * 640 + col) <= 265936) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265937 && (row * 640 + col) <= 265951) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 265952 && (row * 640 + col) <= 265952) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265953 && (row * 640 + col) <= 265962) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 265963 && (row * 640 + col) <= 265963) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265964 && (row * 640 + col) <= 265980) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 265981 && (row * 640 + col) <= 265981) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 265982 && (row * 640 + col) <= 266575) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 266576 && (row * 640 + col) <= 266576) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 266577 && (row * 640 + col) <= 266591) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 266592 && (row * 640 + col) <= 266592) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 266593 && (row * 640 + col) <= 266602) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 266603 && (row * 640 + col) <= 266603) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 266604 && (row * 640 + col) <= 266620) color_data <= 12'b101101110101; else
        if ((row * 640 + col) >= 266621 && (row * 640 + col) <= 266621) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 266622 && (row * 640 + col) <= 267215) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 267216 && (row * 640 + col) <= 267232) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 267233 && (row * 640 + col) <= 267242) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 267243 && (row * 640 + col) <= 267261) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 267262 && (row * 640 + col) <= 284159) color_data <= 12'b101010101010; else
        if ((row * 640 + col) >= 284160 && (row * 640 + col) < 307200) color_data <= 12'b010010000001; else
        color_data <= 12'b000000000000;
    end
endmodule
