module game_over_rom (
	input wire clk,
    input wire [7:0] row,
    input wire [8:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 346 + col) >= 0 && (row * 346 + col) <= 362) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 675 && (row * 346 + col) <= 708) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 1021 && (row * 346 + col) <= 1054) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 1057 && (row * 346 + col) <= 1364) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 1367 && (row * 346 + col) <= 1400) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 1403 && (row * 346 + col) <= 1710) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 1713 && (row * 346 + col) <= 1738) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 1749 && (row * 346 + col) <= 2056) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 2067 && (row * 346 + col) <= 2084) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 2095 && (row * 346 + col) <= 2402) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 2413 && (row * 346 + col) <= 2430) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 2433 && (row * 346 + col) <= 2756) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 2759 && (row * 346 + col) <= 2776) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 2779 && (row * 346 + col) <= 3102) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 3105 && (row * 346 + col) <= 3118) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 3125 && (row * 346 + col) <= 3448) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 3455 && (row * 346 + col) <= 3464) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 3471 && (row * 346 + col) <= 3794) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 3801 && (row * 346 + col) <= 3810) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 3813 && (row * 346 + col) <= 4144) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 4147 && (row * 346 + col) <= 4156) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 4159 && (row * 346 + col) <= 4490) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 4493 && (row * 346 + col) <= 4502) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 4505 && (row * 346 + col) <= 4836) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 4839 && (row * 346 + col) <= 4848) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 4851 && (row * 346 + col) <= 5182) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 5185 && (row * 346 + col) <= 5194) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 5197 && (row * 346 + col) <= 5528) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 5531 && (row * 346 + col) <= 5540) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 5543 && (row * 346 + col) <= 5874) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 5877 && (row * 346 + col) <= 5882) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 5889 && (row * 346 + col) <= 6220) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 6227 && (row * 346 + col) <= 6228) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 6235 && (row * 346 + col) <= 6566) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 6573 && (row * 346 + col) <= 6574) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 6577 && (row * 346 + col) <= 6916) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 6919 && (row * 346 + col) <= 6920) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 6923 && (row * 346 + col) <= 7262) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 7265 && (row * 346 + col) <= 7266) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 7269 && (row * 346 + col) <= 7608) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 7611 && (row * 346 + col) <= 7612) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 7615 && (row * 346 + col) <= 7954) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 7957 && (row * 346 + col) <= 7958) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 7961 && (row * 346 + col) <= 8300) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 8303 && (row * 346 + col) <= 8304) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 8307 && (row * 346 + col) <= 8646) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 8649 && (row * 346 + col) <= 8650) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 8653 && (row * 346 + col) <= 8992) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 8995 && (row * 346 + col) <= 8996) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 8999 && (row * 346 + col) <= 9338) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9341 && (row * 346 + col) <= 9342) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 9345 && (row * 346 + col) <= 9684) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9687 && (row * 346 + col) <= 9688) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 9691 && (row * 346 + col) <= 9706) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9737 && (row * 346 + col) <= 9742) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9773 && (row * 346 + col) <= 9778) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9791 && (row * 346 + col) <= 9808) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9821 && (row * 346 + col) <= 9826) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9857 && (row * 346 + col) <= 9874) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9905 && (row * 346 + col) <= 9910) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9923 && (row * 346 + col) <= 9928) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9941 && (row * 346 + col) <= 9946) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 9977 && (row * 346 + col) <= 9982) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10013 && (row * 346 + col) <= 10030) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10033 && (row * 346 + col) <= 10034) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 10037 && (row * 346 + col) <= 10052) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10083 && (row * 346 + col) <= 10088) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10119 && (row * 346 + col) <= 10124) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10137 && (row * 346 + col) <= 10154) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10167 && (row * 346 + col) <= 10172) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10203 && (row * 346 + col) <= 10220) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10251 && (row * 346 + col) <= 10256) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10269 && (row * 346 + col) <= 10274) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10287 && (row * 346 + col) <= 10292) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10323 && (row * 346 + col) <= 10328) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10359 && (row * 346 + col) <= 10376) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10379 && (row * 346 + col) <= 10380) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 10383 && (row * 346 + col) <= 10398) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10429 && (row * 346 + col) <= 10434) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10465 && (row * 346 + col) <= 10470) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10483 && (row * 346 + col) <= 10500) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10513 && (row * 346 + col) <= 10518) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10549 && (row * 346 + col) <= 10566) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10597 && (row * 346 + col) <= 10602) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10615 && (row * 346 + col) <= 10620) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10633 && (row * 346 + col) <= 10638) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10669 && (row * 346 + col) <= 10674) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10705 && (row * 346 + col) <= 10722) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10725 && (row * 346 + col) <= 10726) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 10729 && (row * 346 + col) <= 10744) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10775 && (row * 346 + col) <= 10780) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10811 && (row * 346 + col) <= 10816) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10829 && (row * 346 + col) <= 10846) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10859 && (row * 346 + col) <= 10864) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10895 && (row * 346 + col) <= 10912) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10943 && (row * 346 + col) <= 10948) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10961 && (row * 346 + col) <= 10966) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 10979 && (row * 346 + col) <= 10984) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11015 && (row * 346 + col) <= 11020) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11051 && (row * 346 + col) <= 11068) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11071 && (row * 346 + col) <= 11072) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 11075 && (row * 346 + col) <= 11090) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11121 && (row * 346 + col) <= 11126) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11157 && (row * 346 + col) <= 11162) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11175 && (row * 346 + col) <= 11192) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11205 && (row * 346 + col) <= 11210) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11241 && (row * 346 + col) <= 11258) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11289 && (row * 346 + col) <= 11294) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11307 && (row * 346 + col) <= 11312) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11325 && (row * 346 + col) <= 11330) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11361 && (row * 346 + col) <= 11366) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11397 && (row * 346 + col) <= 11414) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11417 && (row * 346 + col) <= 11418) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 11421 && (row * 346 + col) <= 11436) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11467 && (row * 346 + col) <= 11472) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11503 && (row * 346 + col) <= 11508) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11521 && (row * 346 + col) <= 11538) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11551 && (row * 346 + col) <= 11556) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11587 && (row * 346 + col) <= 11604) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11635 && (row * 346 + col) <= 11640) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11653 && (row * 346 + col) <= 11658) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11671 && (row * 346 + col) <= 11676) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11707 && (row * 346 + col) <= 11712) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11743 && (row * 346 + col) <= 11760) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11763 && (row * 346 + col) <= 11764) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 11767 && (row * 346 + col) <= 11782) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11795 && (row * 346 + col) <= 11800) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11813 && (row * 346 + col) <= 11818) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11831 && (row * 346 + col) <= 11836) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11849 && (row * 346 + col) <= 11854) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11873 && (row * 346 + col) <= 11878) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11897 && (row * 346 + col) <= 11902) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11915 && (row * 346 + col) <= 11920) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11933 && (row * 346 + col) <= 11950) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11963 && (row * 346 + col) <= 11968) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11981 && (row * 346 + col) <= 11986) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 11999 && (row * 346 + col) <= 12004) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12017 && (row * 346 + col) <= 12022) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12035 && (row * 346 + col) <= 12040) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12053 && (row * 346 + col) <= 12058) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12071 && (row * 346 + col) <= 12076) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12089 && (row * 346 + col) <= 12106) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12109 && (row * 346 + col) <= 12110) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 12113 && (row * 346 + col) <= 12128) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12141 && (row * 346 + col) <= 12146) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12159 && (row * 346 + col) <= 12164) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12177 && (row * 346 + col) <= 12182) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12195 && (row * 346 + col) <= 12200) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12219 && (row * 346 + col) <= 12224) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12243 && (row * 346 + col) <= 12248) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12261 && (row * 346 + col) <= 12266) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12279 && (row * 346 + col) <= 12296) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12309 && (row * 346 + col) <= 12314) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12327 && (row * 346 + col) <= 12332) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12345 && (row * 346 + col) <= 12350) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12363 && (row * 346 + col) <= 12368) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12381 && (row * 346 + col) <= 12386) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12399 && (row * 346 + col) <= 12404) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12417 && (row * 346 + col) <= 12422) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12435 && (row * 346 + col) <= 12452) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12455 && (row * 346 + col) <= 12456) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 12459 && (row * 346 + col) <= 12474) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12487 && (row * 346 + col) <= 12492) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12505 && (row * 346 + col) <= 12510) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12523 && (row * 346 + col) <= 12528) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12541 && (row * 346 + col) <= 12546) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12565 && (row * 346 + col) <= 12570) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12589 && (row * 346 + col) <= 12594) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12607 && (row * 346 + col) <= 12612) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12625 && (row * 346 + col) <= 12642) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12655 && (row * 346 + col) <= 12660) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12673 && (row * 346 + col) <= 12678) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12691 && (row * 346 + col) <= 12696) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12709 && (row * 346 + col) <= 12714) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12727 && (row * 346 + col) <= 12732) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12745 && (row * 346 + col) <= 12750) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12763 && (row * 346 + col) <= 12768) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12781 && (row * 346 + col) <= 12798) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12801 && (row * 346 + col) <= 12802) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 12805 && (row * 346 + col) <= 12820) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12833 && (row * 346 + col) <= 12838) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12851 && (row * 346 + col) <= 12856) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12869 && (row * 346 + col) <= 12874) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12887 && (row * 346 + col) <= 12892) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12911 && (row * 346 + col) <= 12916) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12935 && (row * 346 + col) <= 12940) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12953 && (row * 346 + col) <= 12958) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 12971 && (row * 346 + col) <= 12988) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13001 && (row * 346 + col) <= 13006) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13019 && (row * 346 + col) <= 13024) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13037 && (row * 346 + col) <= 13042) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13055 && (row * 346 + col) <= 13060) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13073 && (row * 346 + col) <= 13078) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13091 && (row * 346 + col) <= 13096) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13109 && (row * 346 + col) <= 13114) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13127 && (row * 346 + col) <= 13144) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13147 && (row * 346 + col) <= 13148) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 13151 && (row * 346 + col) <= 13166) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13179 && (row * 346 + col) <= 13184) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13197 && (row * 346 + col) <= 13202) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13215 && (row * 346 + col) <= 13220) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13233 && (row * 346 + col) <= 13238) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13257 && (row * 346 + col) <= 13262) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13281 && (row * 346 + col) <= 13286) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13299 && (row * 346 + col) <= 13304) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13317 && (row * 346 + col) <= 13334) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13347 && (row * 346 + col) <= 13352) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13365 && (row * 346 + col) <= 13370) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13383 && (row * 346 + col) <= 13388) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13401 && (row * 346 + col) <= 13406) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13419 && (row * 346 + col) <= 13424) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13437 && (row * 346 + col) <= 13442) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13455 && (row * 346 + col) <= 13460) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13473 && (row * 346 + col) <= 13490) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13493 && (row * 346 + col) <= 13494) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 13497 && (row * 346 + col) <= 13512) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13525 && (row * 346 + col) <= 13530) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13543 && (row * 346 + col) <= 13548) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13561 && (row * 346 + col) <= 13566) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13579 && (row * 346 + col) <= 13584) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13603 && (row * 346 + col) <= 13608) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13627 && (row * 346 + col) <= 13632) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13645 && (row * 346 + col) <= 13650) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13663 && (row * 346 + col) <= 13680) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13693 && (row * 346 + col) <= 13698) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13711 && (row * 346 + col) <= 13716) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13729 && (row * 346 + col) <= 13734) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13747 && (row * 346 + col) <= 13752) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13765 && (row * 346 + col) <= 13770) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13783 && (row * 346 + col) <= 13788) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13801 && (row * 346 + col) <= 13806) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13819 && (row * 346 + col) <= 13836) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13839 && (row * 346 + col) <= 13840) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 13843 && (row * 346 + col) <= 13858) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13871 && (row * 346 + col) <= 13894) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13907 && (row * 346 + col) <= 13912) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13925 && (row * 346 + col) <= 13930) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13973 && (row * 346 + col) <= 13978) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 13991 && (row * 346 + col) <= 14026) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14039 && (row * 346 + col) <= 14044) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14057 && (row * 346 + col) <= 14062) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14075 && (row * 346 + col) <= 14080) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14093 && (row * 346 + col) <= 14098) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14111 && (row * 346 + col) <= 14134) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14147 && (row * 346 + col) <= 14152) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14165 && (row * 346 + col) <= 14182) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14185 && (row * 346 + col) <= 14186) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 14189 && (row * 346 + col) <= 14204) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14217 && (row * 346 + col) <= 14240) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14253 && (row * 346 + col) <= 14258) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14271 && (row * 346 + col) <= 14276) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14319 && (row * 346 + col) <= 14324) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14337 && (row * 346 + col) <= 14372) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14385 && (row * 346 + col) <= 14390) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14403 && (row * 346 + col) <= 14408) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14421 && (row * 346 + col) <= 14426) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14439 && (row * 346 + col) <= 14444) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14457 && (row * 346 + col) <= 14480) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14493 && (row * 346 + col) <= 14498) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14511 && (row * 346 + col) <= 14528) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14531 && (row * 346 + col) <= 14532) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 14535 && (row * 346 + col) <= 14550) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14563 && (row * 346 + col) <= 14586) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14599 && (row * 346 + col) <= 14604) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14617 && (row * 346 + col) <= 14622) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14665 && (row * 346 + col) <= 14670) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14683 && (row * 346 + col) <= 14718) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14731 && (row * 346 + col) <= 14736) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14749 && (row * 346 + col) <= 14754) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14767 && (row * 346 + col) <= 14772) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14785 && (row * 346 + col) <= 14790) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14803 && (row * 346 + col) <= 14826) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14839 && (row * 346 + col) <= 14844) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14857 && (row * 346 + col) <= 14874) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14877 && (row * 346 + col) <= 14878) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 14881 && (row * 346 + col) <= 14896) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14909 && (row * 346 + col) <= 14932) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14945 && (row * 346 + col) <= 14950) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 14963 && (row * 346 + col) <= 14968) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15011 && (row * 346 + col) <= 15016) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15029 && (row * 346 + col) <= 15064) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15077 && (row * 346 + col) <= 15082) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15095 && (row * 346 + col) <= 15100) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15113 && (row * 346 + col) <= 15118) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15131 && (row * 346 + col) <= 15136) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15149 && (row * 346 + col) <= 15172) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15185 && (row * 346 + col) <= 15190) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15203 && (row * 346 + col) <= 15220) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15223 && (row * 346 + col) <= 15224) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 15227 && (row * 346 + col) <= 15242) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15255 && (row * 346 + col) <= 15278) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15291 && (row * 346 + col) <= 15296) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15309 && (row * 346 + col) <= 15314) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15357 && (row * 346 + col) <= 15362) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15375 && (row * 346 + col) <= 15410) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15423 && (row * 346 + col) <= 15428) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15441 && (row * 346 + col) <= 15446) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15459 && (row * 346 + col) <= 15464) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15477 && (row * 346 + col) <= 15482) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15495 && (row * 346 + col) <= 15518) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15531 && (row * 346 + col) <= 15536) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15549 && (row * 346 + col) <= 15566) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15569 && (row * 346 + col) <= 15570) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 15573 && (row * 346 + col) <= 15588) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15601 && (row * 346 + col) <= 15624) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15637 && (row * 346 + col) <= 15642) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15655 && (row * 346 + col) <= 15660) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15703 && (row * 346 + col) <= 15708) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15721 && (row * 346 + col) <= 15756) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15769 && (row * 346 + col) <= 15774) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15787 && (row * 346 + col) <= 15792) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15805 && (row * 346 + col) <= 15810) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15823 && (row * 346 + col) <= 15828) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15841 && (row * 346 + col) <= 15864) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15877 && (row * 346 + col) <= 15882) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15895 && (row * 346 + col) <= 15912) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15915 && (row * 346 + col) <= 15916) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 15919 && (row * 346 + col) <= 15934) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15947 && (row * 346 + col) <= 15950) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 15965 && (row * 346 + col) <= 15970) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16001 && (row * 346 + col) <= 16006) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16019 && (row * 346 + col) <= 16024) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16031 && (row * 346 + col) <= 16036) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16049 && (row * 346 + col) <= 16054) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16079 && (row * 346 + col) <= 16102) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16115 && (row * 346 + col) <= 16120) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16133 && (row * 346 + col) <= 16138) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16151 && (row * 346 + col) <= 16156) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16169 && (row * 346 + col) <= 16174) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16199 && (row * 346 + col) <= 16210) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16235 && (row * 346 + col) <= 16258) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16261 && (row * 346 + col) <= 16262) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 16265 && (row * 346 + col) <= 16280) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16293 && (row * 346 + col) <= 16296) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16311 && (row * 346 + col) <= 16316) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16347 && (row * 346 + col) <= 16352) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16365 && (row * 346 + col) <= 16370) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16377 && (row * 346 + col) <= 16382) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16395 && (row * 346 + col) <= 16400) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16425 && (row * 346 + col) <= 16448) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16461 && (row * 346 + col) <= 16466) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16479 && (row * 346 + col) <= 16484) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16497 && (row * 346 + col) <= 16502) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16515 && (row * 346 + col) <= 16520) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16545 && (row * 346 + col) <= 16556) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16581 && (row * 346 + col) <= 16604) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16607 && (row * 346 + col) <= 16608) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 16611 && (row * 346 + col) <= 16626) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16639 && (row * 346 + col) <= 16642) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16657 && (row * 346 + col) <= 16662) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16693 && (row * 346 + col) <= 16698) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16711 && (row * 346 + col) <= 16716) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16723 && (row * 346 + col) <= 16728) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16741 && (row * 346 + col) <= 16746) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16771 && (row * 346 + col) <= 16794) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16807 && (row * 346 + col) <= 16812) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16825 && (row * 346 + col) <= 16830) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16843 && (row * 346 + col) <= 16848) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16861 && (row * 346 + col) <= 16866) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16891 && (row * 346 + col) <= 16902) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16927 && (row * 346 + col) <= 16950) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16953 && (row * 346 + col) <= 16954) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 16957 && (row * 346 + col) <= 16972) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 16985 && (row * 346 + col) <= 16988) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17003 && (row * 346 + col) <= 17008) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17039 && (row * 346 + col) <= 17044) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17057 && (row * 346 + col) <= 17062) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17069 && (row * 346 + col) <= 17074) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17087 && (row * 346 + col) <= 17092) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17117 && (row * 346 + col) <= 17140) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17153 && (row * 346 + col) <= 17158) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17171 && (row * 346 + col) <= 17176) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17189 && (row * 346 + col) <= 17194) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17207 && (row * 346 + col) <= 17212) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17237 && (row * 346 + col) <= 17248) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17273 && (row * 346 + col) <= 17296) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17299 && (row * 346 + col) <= 17300) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 17303 && (row * 346 + col) <= 17318) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17331 && (row * 346 + col) <= 17334) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17349 && (row * 346 + col) <= 17354) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17385 && (row * 346 + col) <= 17390) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17403 && (row * 346 + col) <= 17408) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17415 && (row * 346 + col) <= 17420) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17433 && (row * 346 + col) <= 17438) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17463 && (row * 346 + col) <= 17486) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17499 && (row * 346 + col) <= 17504) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17517 && (row * 346 + col) <= 17522) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17535 && (row * 346 + col) <= 17540) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17553 && (row * 346 + col) <= 17558) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17583 && (row * 346 + col) <= 17594) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17619 && (row * 346 + col) <= 17642) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17645 && (row * 346 + col) <= 17646) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 17649 && (row * 346 + col) <= 17664) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17677 && (row * 346 + col) <= 17680) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17695 && (row * 346 + col) <= 17700) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17731 && (row * 346 + col) <= 17736) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17749 && (row * 346 + col) <= 17754) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17761 && (row * 346 + col) <= 17766) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17779 && (row * 346 + col) <= 17784) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17809 && (row * 346 + col) <= 17832) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17845 && (row * 346 + col) <= 17850) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17863 && (row * 346 + col) <= 17868) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17881 && (row * 346 + col) <= 17886) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17899 && (row * 346 + col) <= 17904) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17929 && (row * 346 + col) <= 17940) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17965 && (row * 346 + col) <= 17988) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 17991 && (row * 346 + col) <= 17992) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 17995 && (row * 346 + col) <= 18010) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18023 && (row * 346 + col) <= 18028) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18041 && (row * 346 + col) <= 18046) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18059 && (row * 346 + col) <= 18064) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18077 && (row * 346 + col) <= 18082) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18095 && (row * 346 + col) <= 18112) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18125 && (row * 346 + col) <= 18130) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18143 && (row * 346 + col) <= 18178) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18191 && (row * 346 + col) <= 18196) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18209 && (row * 346 + col) <= 18214) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18227 && (row * 346 + col) <= 18232) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18245 && (row * 346 + col) <= 18250) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18263 && (row * 346 + col) <= 18286) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18299 && (row * 346 + col) <= 18304) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18317 && (row * 346 + col) <= 18334) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18337 && (row * 346 + col) <= 18338) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 18341 && (row * 346 + col) <= 18356) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18369 && (row * 346 + col) <= 18374) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18387 && (row * 346 + col) <= 18392) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18405 && (row * 346 + col) <= 18410) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18423 && (row * 346 + col) <= 18428) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18441 && (row * 346 + col) <= 18458) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18471 && (row * 346 + col) <= 18476) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18489 && (row * 346 + col) <= 18524) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18537 && (row * 346 + col) <= 18542) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18555 && (row * 346 + col) <= 18560) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18573 && (row * 346 + col) <= 18578) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18591 && (row * 346 + col) <= 18596) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18609 && (row * 346 + col) <= 18632) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18645 && (row * 346 + col) <= 18650) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18663 && (row * 346 + col) <= 18680) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18683 && (row * 346 + col) <= 18684) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 18687 && (row * 346 + col) <= 18702) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18715 && (row * 346 + col) <= 18720) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18733 && (row * 346 + col) <= 18738) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18751 && (row * 346 + col) <= 18756) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18769 && (row * 346 + col) <= 18774) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18787 && (row * 346 + col) <= 18804) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18817 && (row * 346 + col) <= 18822) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18835 && (row * 346 + col) <= 18870) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18883 && (row * 346 + col) <= 18888) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18901 && (row * 346 + col) <= 18906) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18919 && (row * 346 + col) <= 18924) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18937 && (row * 346 + col) <= 18942) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18955 && (row * 346 + col) <= 18978) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 18991 && (row * 346 + col) <= 18996) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19009 && (row * 346 + col) <= 19026) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19029 && (row * 346 + col) <= 19030) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 19033 && (row * 346 + col) <= 19048) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19061 && (row * 346 + col) <= 19066) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19079 && (row * 346 + col) <= 19084) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19097 && (row * 346 + col) <= 19102) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19115 && (row * 346 + col) <= 19120) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19133 && (row * 346 + col) <= 19150) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19163 && (row * 346 + col) <= 19168) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19181 && (row * 346 + col) <= 19216) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19229 && (row * 346 + col) <= 19234) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19247 && (row * 346 + col) <= 19252) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19265 && (row * 346 + col) <= 19270) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19283 && (row * 346 + col) <= 19288) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19301 && (row * 346 + col) <= 19324) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19337 && (row * 346 + col) <= 19342) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19355 && (row * 346 + col) <= 19372) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19375 && (row * 346 + col) <= 19376) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 19379 && (row * 346 + col) <= 19394) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19407 && (row * 346 + col) <= 19412) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19425 && (row * 346 + col) <= 19430) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19443 && (row * 346 + col) <= 19448) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19461 && (row * 346 + col) <= 19466) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19479 && (row * 346 + col) <= 19496) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19509 && (row * 346 + col) <= 19514) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19527 && (row * 346 + col) <= 19562) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19575 && (row * 346 + col) <= 19580) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19593 && (row * 346 + col) <= 19598) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19611 && (row * 346 + col) <= 19616) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19629 && (row * 346 + col) <= 19634) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19647 && (row * 346 + col) <= 19670) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19683 && (row * 346 + col) <= 19688) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19701 && (row * 346 + col) <= 19718) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19721 && (row * 346 + col) <= 19722) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 19725 && (row * 346 + col) <= 19740) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19753 && (row * 346 + col) <= 19758) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19771 && (row * 346 + col) <= 19776) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19789 && (row * 346 + col) <= 19794) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19807 && (row * 346 + col) <= 19812) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19825 && (row * 346 + col) <= 19842) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19855 && (row * 346 + col) <= 19860) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19873 && (row * 346 + col) <= 19908) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19921 && (row * 346 + col) <= 19926) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19939 && (row * 346 + col) <= 19944) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19957 && (row * 346 + col) <= 19962) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19975 && (row * 346 + col) <= 19980) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 19993 && (row * 346 + col) <= 20016) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20029 && (row * 346 + col) <= 20034) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20047 && (row * 346 + col) <= 20064) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20067 && (row * 346 + col) <= 20068) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 20071 && (row * 346 + col) <= 20086) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20099 && (row * 346 + col) <= 20104) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20117 && (row * 346 + col) <= 20122) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20135 && (row * 346 + col) <= 20140) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20153 && (row * 346 + col) <= 20158) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20171 && (row * 346 + col) <= 20188) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20201 && (row * 346 + col) <= 20206) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20219 && (row * 346 + col) <= 20254) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20267 && (row * 346 + col) <= 20272) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20285 && (row * 346 + col) <= 20290) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20303 && (row * 346 + col) <= 20308) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20321 && (row * 346 + col) <= 20326) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20339 && (row * 346 + col) <= 20362) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20375 && (row * 346 + col) <= 20380) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20393 && (row * 346 + col) <= 20410) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20413 && (row * 346 + col) <= 20414) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 20417 && (row * 346 + col) <= 20432) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20445 && (row * 346 + col) <= 20450) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20463 && (row * 346 + col) <= 20468) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20481 && (row * 346 + col) <= 20486) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20499 && (row * 346 + col) <= 20504) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20517 && (row * 346 + col) <= 20534) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20547 && (row * 346 + col) <= 20552) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20565 && (row * 346 + col) <= 20600) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20613 && (row * 346 + col) <= 20618) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20631 && (row * 346 + col) <= 20636) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20649 && (row * 346 + col) <= 20654) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20667 && (row * 346 + col) <= 20672) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20685 && (row * 346 + col) <= 20708) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20721 && (row * 346 + col) <= 20726) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20739 && (row * 346 + col) <= 20756) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20759 && (row * 346 + col) <= 20760) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 20763 && (row * 346 + col) <= 20778) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20791 && (row * 346 + col) <= 20796) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20809 && (row * 346 + col) <= 20814) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20827 && (row * 346 + col) <= 20832) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20845 && (row * 346 + col) <= 20850) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20863 && (row * 346 + col) <= 20880) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20893 && (row * 346 + col) <= 20898) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20911 && (row * 346 + col) <= 20946) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20959 && (row * 346 + col) <= 20964) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20977 && (row * 346 + col) <= 20982) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 20995 && (row * 346 + col) <= 21000) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21013 && (row * 346 + col) <= 21018) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21031 && (row * 346 + col) <= 21054) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21067 && (row * 346 + col) <= 21072) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21085 && (row * 346 + col) <= 21102) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21105 && (row * 346 + col) <= 21106) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 21109 && (row * 346 + col) <= 21124) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21137 && (row * 346 + col) <= 21142) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21155 && (row * 346 + col) <= 21160) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21173 && (row * 346 + col) <= 21178) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21191 && (row * 346 + col) <= 21196) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21209 && (row * 346 + col) <= 21226) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21239 && (row * 346 + col) <= 21244) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21257 && (row * 346 + col) <= 21292) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21305 && (row * 346 + col) <= 21310) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21323 && (row * 346 + col) <= 21328) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21341 && (row * 346 + col) <= 21346) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21359 && (row * 346 + col) <= 21364) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21377 && (row * 346 + col) <= 21400) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21413 && (row * 346 + col) <= 21418) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21431 && (row * 346 + col) <= 21448) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21451 && (row * 346 + col) <= 21452) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 21455 && (row * 346 + col) <= 21470) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21483 && (row * 346 + col) <= 21488) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21501 && (row * 346 + col) <= 21506) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21519 && (row * 346 + col) <= 21524) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21537 && (row * 346 + col) <= 21542) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21555 && (row * 346 + col) <= 21572) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21585 && (row * 346 + col) <= 21590) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21603 && (row * 346 + col) <= 21638) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21651 && (row * 346 + col) <= 21656) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21669 && (row * 346 + col) <= 21674) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21687 && (row * 346 + col) <= 21692) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21705 && (row * 346 + col) <= 21710) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21723 && (row * 346 + col) <= 21746) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21759 && (row * 346 + col) <= 21764) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21777 && (row * 346 + col) <= 21794) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21797 && (row * 346 + col) <= 21798) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 21801 && (row * 346 + col) <= 21816) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21829 && (row * 346 + col) <= 21834) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21847 && (row * 346 + col) <= 21852) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21865 && (row * 346 + col) <= 21870) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21883 && (row * 346 + col) <= 21888) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21901 && (row * 346 + col) <= 21918) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21931 && (row * 346 + col) <= 21936) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21949 && (row * 346 + col) <= 21984) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 21997 && (row * 346 + col) <= 22002) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22015 && (row * 346 + col) <= 22020) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22033 && (row * 346 + col) <= 22038) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22051 && (row * 346 + col) <= 22056) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22069 && (row * 346 + col) <= 22092) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22105 && (row * 346 + col) <= 22110) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22123 && (row * 346 + col) <= 22140) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22143 && (row * 346 + col) <= 22144) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 22147 && (row * 346 + col) <= 22162) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22175 && (row * 346 + col) <= 22180) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22193 && (row * 346 + col) <= 22198) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22211 && (row * 346 + col) <= 22216) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22229 && (row * 346 + col) <= 22234) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22247 && (row * 346 + col) <= 22264) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22277 && (row * 346 + col) <= 22282) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22295 && (row * 346 + col) <= 22300) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22313 && (row * 346 + col) <= 22330) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22343 && (row * 346 + col) <= 22348) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22361 && (row * 346 + col) <= 22372) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22391 && (row * 346 + col) <= 22402) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22415 && (row * 346 + col) <= 22420) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22433 && (row * 346 + col) <= 22438) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22451 && (row * 346 + col) <= 22456) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22469 && (row * 346 + col) <= 22486) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22489 && (row * 346 + col) <= 22490) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 22493 && (row * 346 + col) <= 22508) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22521 && (row * 346 + col) <= 22526) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22539 && (row * 346 + col) <= 22544) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22557 && (row * 346 + col) <= 22562) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22575 && (row * 346 + col) <= 22580) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22593 && (row * 346 + col) <= 22610) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22623 && (row * 346 + col) <= 22628) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22641 && (row * 346 + col) <= 22646) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22659 && (row * 346 + col) <= 22676) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22689 && (row * 346 + col) <= 22694) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22707 && (row * 346 + col) <= 22718) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22737 && (row * 346 + col) <= 22748) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22761 && (row * 346 + col) <= 22766) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22779 && (row * 346 + col) <= 22784) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22797 && (row * 346 + col) <= 22802) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22815 && (row * 346 + col) <= 22832) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22835 && (row * 346 + col) <= 22836) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 22839 && (row * 346 + col) <= 22854) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22867 && (row * 346 + col) <= 22872) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22885 && (row * 346 + col) <= 22890) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22903 && (row * 346 + col) <= 22908) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22921 && (row * 346 + col) <= 22926) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22939 && (row * 346 + col) <= 22956) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22969 && (row * 346 + col) <= 22974) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 22987 && (row * 346 + col) <= 22992) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23005 && (row * 346 + col) <= 23022) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23035 && (row * 346 + col) <= 23040) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23053 && (row * 346 + col) <= 23064) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23083 && (row * 346 + col) <= 23094) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23107 && (row * 346 + col) <= 23112) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23125 && (row * 346 + col) <= 23130) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23143 && (row * 346 + col) <= 23148) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23161 && (row * 346 + col) <= 23178) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23181 && (row * 346 + col) <= 23182) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 23185 && (row * 346 + col) <= 23200) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23213 && (row * 346 + col) <= 23218) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23231 && (row * 346 + col) <= 23236) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23249 && (row * 346 + col) <= 23254) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23267 && (row * 346 + col) <= 23272) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23285 && (row * 346 + col) <= 23302) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23315 && (row * 346 + col) <= 23320) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23333 && (row * 346 + col) <= 23338) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23351 && (row * 346 + col) <= 23368) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23381 && (row * 346 + col) <= 23386) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23399 && (row * 346 + col) <= 23410) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23429 && (row * 346 + col) <= 23440) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23453 && (row * 346 + col) <= 23458) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23471 && (row * 346 + col) <= 23476) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23489 && (row * 346 + col) <= 23494) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23507 && (row * 346 + col) <= 23524) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23527 && (row * 346 + col) <= 23528) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 23531 && (row * 346 + col) <= 23546) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23559 && (row * 346 + col) <= 23564) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23577 && (row * 346 + col) <= 23582) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23595 && (row * 346 + col) <= 23600) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23613 && (row * 346 + col) <= 23618) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23631 && (row * 346 + col) <= 23648) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23661 && (row * 346 + col) <= 23666) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23679 && (row * 346 + col) <= 23684) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23697 && (row * 346 + col) <= 23714) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23727 && (row * 346 + col) <= 23732) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23745 && (row * 346 + col) <= 23756) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23775 && (row * 346 + col) <= 23786) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23799 && (row * 346 + col) <= 23804) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23817 && (row * 346 + col) <= 23822) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23835 && (row * 346 + col) <= 23840) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23853 && (row * 346 + col) <= 23870) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23873 && (row * 346 + col) <= 23874) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 23877 && (row * 346 + col) <= 23892) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23905 && (row * 346 + col) <= 23910) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23923 && (row * 346 + col) <= 23928) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23941 && (row * 346 + col) <= 23946) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23959 && (row * 346 + col) <= 23964) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 23977 && (row * 346 + col) <= 23994) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24007 && (row * 346 + col) <= 24012) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24025 && (row * 346 + col) <= 24030) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24043 && (row * 346 + col) <= 24060) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24073 && (row * 346 + col) <= 24078) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24091 && (row * 346 + col) <= 24102) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24121 && (row * 346 + col) <= 24132) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24145 && (row * 346 + col) <= 24150) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24163 && (row * 346 + col) <= 24168) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24181 && (row * 346 + col) <= 24186) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24199 && (row * 346 + col) <= 24216) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24219 && (row * 346 + col) <= 24220) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 24223 && (row * 346 + col) <= 24238) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24269 && (row * 346 + col) <= 24274) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24287 && (row * 346 + col) <= 24292) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24305 && (row * 346 + col) <= 24310) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24323 && (row * 346 + col) <= 24340) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24353 && (row * 346 + col) <= 24358) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24389 && (row * 346 + col) <= 24406) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24437 && (row * 346 + col) <= 24448) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24467 && (row * 346 + col) <= 24478) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24509 && (row * 346 + col) <= 24514) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24527 && (row * 346 + col) <= 24532) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24545 && (row * 346 + col) <= 24562) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24565 && (row * 346 + col) <= 24566) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 24569 && (row * 346 + col) <= 24584) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24615 && (row * 346 + col) <= 24620) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24633 && (row * 346 + col) <= 24638) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24651 && (row * 346 + col) <= 24656) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24669 && (row * 346 + col) <= 24686) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24699 && (row * 346 + col) <= 24704) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24735 && (row * 346 + col) <= 24752) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24783 && (row * 346 + col) <= 24794) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24813 && (row * 346 + col) <= 24824) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24855 && (row * 346 + col) <= 24860) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24873 && (row * 346 + col) <= 24878) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24891 && (row * 346 + col) <= 24908) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24911 && (row * 346 + col) <= 24912) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 24915 && (row * 346 + col) <= 24930) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24961 && (row * 346 + col) <= 24966) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24979 && (row * 346 + col) <= 24984) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 24997 && (row * 346 + col) <= 25002) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25015 && (row * 346 + col) <= 25032) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25045 && (row * 346 + col) <= 25050) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25081 && (row * 346 + col) <= 25098) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25129 && (row * 346 + col) <= 25144) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25155 && (row * 346 + col) <= 25170) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25201 && (row * 346 + col) <= 25206) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25219 && (row * 346 + col) <= 25224) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25237 && (row * 346 + col) <= 25254) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25257 && (row * 346 + col) <= 25258) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 25261 && (row * 346 + col) <= 25276) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25307 && (row * 346 + col) <= 25312) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25325 && (row * 346 + col) <= 25330) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25343 && (row * 346 + col) <= 25348) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25361 && (row * 346 + col) <= 25378) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25391 && (row * 346 + col) <= 25396) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25427 && (row * 346 + col) <= 25444) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25475 && (row * 346 + col) <= 25490) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25501 && (row * 346 + col) <= 25516) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25547 && (row * 346 + col) <= 25552) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25565 && (row * 346 + col) <= 25570) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25583 && (row * 346 + col) <= 25600) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25603 && (row * 346 + col) <= 25604) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 25607 && (row * 346 + col) <= 25622) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25653 && (row * 346 + col) <= 25658) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25671 && (row * 346 + col) <= 25676) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25689 && (row * 346 + col) <= 25694) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25707 && (row * 346 + col) <= 25724) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25737 && (row * 346 + col) <= 25742) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25773 && (row * 346 + col) <= 25790) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25821 && (row * 346 + col) <= 25836) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25847 && (row * 346 + col) <= 25862) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25893 && (row * 346 + col) <= 25898) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25911 && (row * 346 + col) <= 25916) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25929 && (row * 346 + col) <= 25946) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25949 && (row * 346 + col) <= 25950) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 25953 && (row * 346 + col) <= 25968) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 25999 && (row * 346 + col) <= 26004) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26017 && (row * 346 + col) <= 26022) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26035 && (row * 346 + col) <= 26040) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26053 && (row * 346 + col) <= 26070) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26083 && (row * 346 + col) <= 26088) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26119 && (row * 346 + col) <= 26136) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26167 && (row * 346 + col) <= 26182) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26193 && (row * 346 + col) <= 26208) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26239 && (row * 346 + col) <= 26244) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26257 && (row * 346 + col) <= 26262) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26275 && (row * 346 + col) <= 26292) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26295 && (row * 346 + col) <= 26296) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 26299 && (row * 346 + col) <= 26638) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26641 && (row * 346 + col) <= 26642) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 26645 && (row * 346 + col) <= 26984) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 26987 && (row * 346 + col) <= 26988) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 26991 && (row * 346 + col) <= 27330) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 27333 && (row * 346 + col) <= 27334) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 27337 && (row * 346 + col) <= 27676) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 27679 && (row * 346 + col) <= 27680) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 27683 && (row * 346 + col) <= 28022) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 28025 && (row * 346 + col) <= 28026) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 28029 && (row * 346 + col) <= 28368) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 28371 && (row * 346 + col) <= 28372) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 28375 && (row * 346 + col) <= 28714) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 28717 && (row * 346 + col) <= 28718) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 28721 && (row * 346 + col) <= 29060) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 29063 && (row * 346 + col) <= 29064) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 29067 && (row * 346 + col) <= 29406) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 29409 && (row * 346 + col) <= 29410) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 29413 && (row * 346 + col) <= 29752) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 29755 && (row * 346 + col) <= 29756) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 29759 && (row * 346 + col) <= 30098) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 30101 && (row * 346 + col) <= 30102) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 30105 && (row * 346 + col) <= 30444) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 30447 && (row * 346 + col) <= 30448) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 30451 && (row * 346 + col) <= 30790) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 30793 && (row * 346 + col) <= 30794) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 30797 && (row * 346 + col) <= 31136) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 31139 && (row * 346 + col) <= 31140) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 31143 && (row * 346 + col) <= 31482) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 31485 && (row * 346 + col) <= 31486) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 31489 && (row * 346 + col) <= 31828) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 31831 && (row * 346 + col) <= 31832) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 31835 && (row * 346 + col) <= 32174) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 32177 && (row * 346 + col) <= 32178) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 32181 && (row * 346 + col) <= 32520) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 32523 && (row * 346 + col) <= 32524) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 32527 && (row * 346 + col) <= 32866) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 32869 && (row * 346 + col) <= 32870) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 32873 && (row * 346 + col) <= 33212) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 33215 && (row * 346 + col) <= 33216) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 33219 && (row * 346 + col) <= 33558) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 33561 && (row * 346 + col) <= 33562) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 33565 && (row * 346 + col) <= 33904) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 33907 && (row * 346 + col) <= 33908) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 33911 && (row * 346 + col) <= 34250) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 34253 && (row * 346 + col) <= 34254) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 34257 && (row * 346 + col) <= 34596) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 34599 && (row * 346 + col) <= 34600) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 34603 && (row * 346 + col) <= 34942) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 34945 && (row * 346 + col) <= 34946) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 34949 && (row * 346 + col) <= 35288) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 35291 && (row * 346 + col) <= 35292) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 35295 && (row * 346 + col) <= 35332) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 35333 && (row * 346 + col) <= 35600) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 35601 && (row * 346 + col) <= 35634) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 35637 && (row * 346 + col) <= 35638) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 35641 && (row * 346 + col) <= 35678) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 35679 && (row * 346 + col) <= 35946) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 35947 && (row * 346 + col) <= 35980) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 35983 && (row * 346 + col) <= 35984) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 35987 && (row * 346 + col) <= 36024) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 36025 && (row * 346 + col) <= 36292) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 36293 && (row * 346 + col) <= 36326) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 36329 && (row * 346 + col) <= 36330) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 36333 && (row * 346 + col) <= 36370) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 36371 && (row * 346 + col) <= 36373) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 36374 && (row * 346 + col) <= 36635) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 36636 && (row * 346 + col) <= 36638) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 36639 && (row * 346 + col) <= 36672) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 36675 && (row * 346 + col) <= 36676) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 36679 && (row * 346 + col) <= 36716) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 36717 && (row * 346 + col) <= 36719) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 36720 && (row * 346 + col) <= 36981) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 36982 && (row * 346 + col) <= 36984) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 36985 && (row * 346 + col) <= 37018) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37021 && (row * 346 + col) <= 37022) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 37025 && (row * 346 + col) <= 37062) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37063 && (row * 346 + col) <= 37065) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 37066 && (row * 346 + col) <= 37327) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37328 && (row * 346 + col) <= 37330) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 37331 && (row * 346 + col) <= 37364) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37367 && (row * 346 + col) <= 37368) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 37371 && (row * 346 + col) <= 37408) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37409 && (row * 346 + col) <= 37411) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 37412 && (row * 346 + col) <= 37673) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37674 && (row * 346 + col) <= 37676) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 37677 && (row * 346 + col) <= 37710) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37713 && (row * 346 + col) <= 37714) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 37717 && (row * 346 + col) <= 37754) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 37755 && (row * 346 + col) <= 37757) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 37758 && (row * 346 + col) <= 38019) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38020 && (row * 346 + col) <= 38022) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 38023 && (row * 346 + col) <= 38056) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38059 && (row * 346 + col) <= 38060) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 38063 && (row * 346 + col) <= 38100) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38101 && (row * 346 + col) <= 38103) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 38104 && (row * 346 + col) <= 38365) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38366 && (row * 346 + col) <= 38368) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 38369 && (row * 346 + col) <= 38402) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38405 && (row * 346 + col) <= 38406) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 38409 && (row * 346 + col) <= 38446) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38447 && (row * 346 + col) <= 38449) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 38450 && (row * 346 + col) <= 38711) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38712 && (row * 346 + col) <= 38714) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 38715 && (row * 346 + col) <= 38748) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38751 && (row * 346 + col) <= 38752) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 38755 && (row * 346 + col) <= 38792) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 38793 && (row * 346 + col) <= 38795) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 38796 && (row * 346 + col) <= 39057) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39058 && (row * 346 + col) <= 39060) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 39061 && (row * 346 + col) <= 39094) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39097 && (row * 346 + col) <= 39098) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 39101 && (row * 346 + col) <= 39138) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39139 && (row * 346 + col) <= 39141) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 39142 && (row * 346 + col) <= 39403) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39404 && (row * 346 + col) <= 39406) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 39407 && (row * 346 + col) <= 39440) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39443 && (row * 346 + col) <= 39444) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 39447 && (row * 346 + col) <= 39484) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39485 && (row * 346 + col) <= 39487) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 39488 && (row * 346 + col) <= 39749) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39750 && (row * 346 + col) <= 39752) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 39753 && (row * 346 + col) <= 39786) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39789 && (row * 346 + col) <= 39790) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 39793 && (row * 346 + col) <= 39830) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 39831 && (row * 346 + col) <= 39833) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 39834 && (row * 346 + col) <= 40095) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40096 && (row * 346 + col) <= 40098) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 40099 && (row * 346 + col) <= 40132) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40135 && (row * 346 + col) <= 40136) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 40139 && (row * 346 + col) <= 40176) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40177 && (row * 346 + col) <= 40179) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 40180 && (row * 346 + col) <= 40204) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40215 && (row * 346 + col) <= 40441) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40442 && (row * 346 + col) <= 40444) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 40445 && (row * 346 + col) <= 40478) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40481 && (row * 346 + col) <= 40482) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 40485 && (row * 346 + col) <= 40522) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40523 && (row * 346 + col) <= 40525) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 40526 && (row * 346 + col) <= 40547) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40564 && (row * 346 + col) <= 40787) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40788 && (row * 346 + col) <= 40790) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 40791 && (row * 346 + col) <= 40824) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40827 && (row * 346 + col) <= 40828) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 40831 && (row * 346 + col) <= 40868) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40869 && (row * 346 + col) <= 40871) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 40872 && (row * 346 + col) <= 40891) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 40898 && (row * 346 + col) <= 40905) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 40912 && (row * 346 + col) <= 41133) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41134 && (row * 346 + col) <= 41136) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41137 && (row * 346 + col) <= 41170) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41173 && (row * 346 + col) <= 41174) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 41177 && (row * 346 + col) <= 41214) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41215 && (row * 346 + col) <= 41217) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41218 && (row * 346 + col) <= 41236) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41241 && (row * 346 + col) <= 41254) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41259 && (row * 346 + col) <= 41479) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41480 && (row * 346 + col) <= 41482) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41483 && (row * 346 + col) <= 41516) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41519 && (row * 346 + col) <= 41520) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 41523 && (row * 346 + col) <= 41560) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41561 && (row * 346 + col) <= 41563) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41564 && (row * 346 + col) <= 41581) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41585 && (row * 346 + col) <= 41602) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41606 && (row * 346 + col) <= 41825) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41826 && (row * 346 + col) <= 41828) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41829 && (row * 346 + col) <= 41862) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41865 && (row * 346 + col) <= 41866) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 41869 && (row * 346 + col) <= 41906) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41907 && (row * 346 + col) <= 41909) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41910 && (row * 346 + col) <= 41926) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 41930 && (row * 346 + col) <= 41949) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 41953 && (row * 346 + col) <= 42171) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42172 && (row * 346 + col) <= 42174) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42175 && (row * 346 + col) <= 42208) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42211 && (row * 346 + col) <= 42212) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 42215 && (row * 346 + col) <= 42252) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42253 && (row * 346 + col) <= 42255) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42256 && (row * 346 + col) <= 42271) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42275 && (row * 346 + col) <= 42296) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42300 && (row * 346 + col) <= 42517) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42518 && (row * 346 + col) <= 42520) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42521 && (row * 346 + col) <= 42554) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42557 && (row * 346 + col) <= 42558) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 42561 && (row * 346 + col) <= 42598) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42599 && (row * 346 + col) <= 42601) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42602 && (row * 346 + col) <= 42616) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42620 && (row * 346 + col) <= 42643) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42647 && (row * 346 + col) <= 42863) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42864 && (row * 346 + col) <= 42866) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42867 && (row * 346 + col) <= 42900) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42903 && (row * 346 + col) <= 42904) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 42907 && (row * 346 + col) <= 42944) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42945 && (row * 346 + col) <= 42947) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42948 && (row * 346 + col) <= 42961) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 42965 && (row * 346 + col) <= 42990) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 42994 && (row * 346 + col) <= 43026) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43042 && (row * 346 + col) <= 43044) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43051 && (row * 346 + col) <= 43062) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43078 && (row * 346 + col) <= 43080) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43087 && (row * 346 + col) <= 43089) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43096 && (row * 346 + col) <= 43110) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43126 && (row * 346 + col) <= 43128) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43144 && (row * 346 + col) <= 43146) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43162 && (row * 346 + col) <= 43164) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43177 && (row * 346 + col) <= 43179) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43186 && (row * 346 + col) <= 43191) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43198 && (row * 346 + col) <= 43209) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43210 && (row * 346 + col) <= 43212) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43213 && (row * 346 + col) <= 43246) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43249 && (row * 346 + col) <= 43250) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 43253 && (row * 346 + col) <= 43290) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43291 && (row * 346 + col) <= 43293) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43294 && (row * 346 + col) <= 43306) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43310 && (row * 346 + col) <= 43337) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43341 && (row * 346 + col) <= 43372) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43388 && (row * 346 + col) <= 43390) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43397 && (row * 346 + col) <= 43408) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43424 && (row * 346 + col) <= 43426) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43433 && (row * 346 + col) <= 43435) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43442 && (row * 346 + col) <= 43456) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43472 && (row * 346 + col) <= 43474) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43490 && (row * 346 + col) <= 43492) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43508 && (row * 346 + col) <= 43510) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43523 && (row * 346 + col) <= 43525) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43532 && (row * 346 + col) <= 43537) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43544 && (row * 346 + col) <= 43555) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43556 && (row * 346 + col) <= 43558) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43559 && (row * 346 + col) <= 43592) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43595 && (row * 346 + col) <= 43596) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 43599 && (row * 346 + col) <= 43636) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43637 && (row * 346 + col) <= 43639) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43640 && (row * 346 + col) <= 43652) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43655 && (row * 346 + col) <= 43684) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43687 && (row * 346 + col) <= 43718) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43734 && (row * 346 + col) <= 43736) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43743 && (row * 346 + col) <= 43754) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43770 && (row * 346 + col) <= 43772) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43779 && (row * 346 + col) <= 43781) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43788 && (row * 346 + col) <= 43802) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43818 && (row * 346 + col) <= 43820) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43836 && (row * 346 + col) <= 43838) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43854 && (row * 346 + col) <= 43856) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43869 && (row * 346 + col) <= 43871) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43878 && (row * 346 + col) <= 43883) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43890 && (row * 346 + col) <= 43901) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43902 && (row * 346 + col) <= 43904) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43905 && (row * 346 + col) <= 43938) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43941 && (row * 346 + col) <= 43942) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 43945 && (row * 346 + col) <= 43982) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 43983 && (row * 346 + col) <= 43985) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 43986 && (row * 346 + col) <= 43997) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44001 && (row * 346 + col) <= 44030) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44034 && (row * 346 + col) <= 44047) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44052 && (row * 346 + col) <= 44064) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44071 && (row * 346 + col) <= 44073) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44080 && (row * 346 + col) <= 44082) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44089 && (row * 346 + col) <= 44100) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44107 && (row * 346 + col) <= 44109) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44116 && (row * 346 + col) <= 44118) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44125 && (row * 346 + col) <= 44127) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44134 && (row * 346 + col) <= 44148) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44155 && (row * 346 + col) <= 44157) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44164 && (row * 346 + col) <= 44166) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44173 && (row * 346 + col) <= 44175) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44182 && (row * 346 + col) <= 44184) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44191 && (row * 346 + col) <= 44193) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44200 && (row * 346 + col) <= 44205) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44212 && (row * 346 + col) <= 44217) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44227 && (row * 346 + col) <= 44229) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44236 && (row * 346 + col) <= 44247) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44248 && (row * 346 + col) <= 44250) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44251 && (row * 346 + col) <= 44284) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44287 && (row * 346 + col) <= 44288) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 44291 && (row * 346 + col) <= 44328) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44329 && (row * 346 + col) <= 44331) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44332 && (row * 346 + col) <= 44343) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44346 && (row * 346 + col) <= 44377) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44380 && (row * 346 + col) <= 44393) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44398 && (row * 346 + col) <= 44410) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44417 && (row * 346 + col) <= 44419) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44426 && (row * 346 + col) <= 44428) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44435 && (row * 346 + col) <= 44446) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44453 && (row * 346 + col) <= 44455) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44462 && (row * 346 + col) <= 44464) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44471 && (row * 346 + col) <= 44473) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44480 && (row * 346 + col) <= 44494) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44501 && (row * 346 + col) <= 44503) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44510 && (row * 346 + col) <= 44512) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44519 && (row * 346 + col) <= 44521) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44528 && (row * 346 + col) <= 44530) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44537 && (row * 346 + col) <= 44539) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44546 && (row * 346 + col) <= 44551) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44558 && (row * 346 + col) <= 44563) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44573 && (row * 346 + col) <= 44575) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44582 && (row * 346 + col) <= 44593) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44594 && (row * 346 + col) <= 44596) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44597 && (row * 346 + col) <= 44630) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44633 && (row * 346 + col) <= 44634) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 44637 && (row * 346 + col) <= 44674) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44675 && (row * 346 + col) <= 44677) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44678 && (row * 346 + col) <= 44689) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44692 && (row * 346 + col) <= 44723) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44726 && (row * 346 + col) <= 44739) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44744 && (row * 346 + col) <= 44756) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44763 && (row * 346 + col) <= 44765) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44772 && (row * 346 + col) <= 44774) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44781 && (row * 346 + col) <= 44792) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44799 && (row * 346 + col) <= 44801) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44808 && (row * 346 + col) <= 44810) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44817 && (row * 346 + col) <= 44819) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44826 && (row * 346 + col) <= 44840) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44847 && (row * 346 + col) <= 44849) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44856 && (row * 346 + col) <= 44858) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44865 && (row * 346 + col) <= 44867) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44874 && (row * 346 + col) <= 44876) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44883 && (row * 346 + col) <= 44885) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44892 && (row * 346 + col) <= 44897) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44904 && (row * 346 + col) <= 44909) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44919 && (row * 346 + col) <= 44921) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44928 && (row * 346 + col) <= 44939) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44940 && (row * 346 + col) <= 44942) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 44943 && (row * 346 + col) <= 44976) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 44979 && (row * 346 + col) <= 44980) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 44983 && (row * 346 + col) <= 45020) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45021 && (row * 346 + col) <= 45023) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45024 && (row * 346 + col) <= 45034) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45038 && (row * 346 + col) <= 45069) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45073 && (row * 346 + col) <= 45085) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45090 && (row * 346 + col) <= 45102) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45109 && (row * 346 + col) <= 45111) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45118 && (row * 346 + col) <= 45120) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45127 && (row * 346 + col) <= 45138) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45145 && (row * 346 + col) <= 45147) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45154 && (row * 346 + col) <= 45156) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45163 && (row * 346 + col) <= 45165) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45172 && (row * 346 + col) <= 45186) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45193 && (row * 346 + col) <= 45195) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45202 && (row * 346 + col) <= 45204) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45211 && (row * 346 + col) <= 45222) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45229 && (row * 346 + col) <= 45231) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45238 && (row * 346 + col) <= 45243) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45250 && (row * 346 + col) <= 45255) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45274 && (row * 346 + col) <= 45285) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45286 && (row * 346 + col) <= 45288) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45289 && (row * 346 + col) <= 45322) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45325 && (row * 346 + col) <= 45326) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 45329 && (row * 346 + col) <= 45366) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45367 && (row * 346 + col) <= 45369) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45370 && (row * 346 + col) <= 45380) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45383 && (row * 346 + col) <= 45386) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45387 && (row * 346 + col) <= 45391) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45392 && (row * 346 + col) <= 45392) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45393 && (row * 346 + col) <= 45396) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45397 && (row * 346 + col) <= 45397) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45398 && (row * 346 + col) <= 45402) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45403 && (row * 346 + col) <= 45403) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45404 && (row * 346 + col) <= 45408) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45409 && (row * 346 + col) <= 45409) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45410 && (row * 346 + col) <= 45413) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45414 && (row * 346 + col) <= 45416) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45419 && (row * 346 + col) <= 45448) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45455 && (row * 346 + col) <= 45457) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45464 && (row * 346 + col) <= 45466) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45473 && (row * 346 + col) <= 45484) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45491 && (row * 346 + col) <= 45493) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45500 && (row * 346 + col) <= 45502) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45509 && (row * 346 + col) <= 45511) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45518 && (row * 346 + col) <= 45532) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45539 && (row * 346 + col) <= 45541) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45548 && (row * 346 + col) <= 45550) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45557 && (row * 346 + col) <= 45568) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45575 && (row * 346 + col) <= 45577) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45584 && (row * 346 + col) <= 45589) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45596 && (row * 346 + col) <= 45601) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45620 && (row * 346 + col) <= 45631) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45632 && (row * 346 + col) <= 45634) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45635 && (row * 346 + col) <= 45668) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45671 && (row * 346 + col) <= 45672) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 45675 && (row * 346 + col) <= 45712) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45713 && (row * 346 + col) <= 45715) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45716 && (row * 346 + col) <= 45726) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45729 && (row * 346 + col) <= 45732) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45733 && (row * 346 + col) <= 45734) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45735 && (row * 346 + col) <= 45735) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45736 && (row * 346 + col) <= 45737) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45738 && (row * 346 + col) <= 45739) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45740 && (row * 346 + col) <= 45741) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45742 && (row * 346 + col) <= 45743) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45744 && (row * 346 + col) <= 45745) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45746 && (row * 346 + col) <= 45746) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45747 && (row * 346 + col) <= 45748) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45749 && (row * 346 + col) <= 45749) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45750 && (row * 346 + col) <= 45751) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45752 && (row * 346 + col) <= 45752) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45753 && (row * 346 + col) <= 45754) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45755 && (row * 346 + col) <= 45756) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45757 && (row * 346 + col) <= 45758) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45759 && (row * 346 + col) <= 45762) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45765 && (row * 346 + col) <= 45794) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45801 && (row * 346 + col) <= 45803) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45810 && (row * 346 + col) <= 45812) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45819 && (row * 346 + col) <= 45830) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45837 && (row * 346 + col) <= 45839) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45846 && (row * 346 + col) <= 45848) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45855 && (row * 346 + col) <= 45857) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45864 && (row * 346 + col) <= 45878) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45885 && (row * 346 + col) <= 45887) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45894 && (row * 346 + col) <= 45896) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45903 && (row * 346 + col) <= 45914) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45921 && (row * 346 + col) <= 45923) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45930 && (row * 346 + col) <= 45935) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45942 && (row * 346 + col) <= 45947) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45966 && (row * 346 + col) <= 45977) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 45978 && (row * 346 + col) <= 45980) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 45981 && (row * 346 + col) <= 46014) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46017 && (row * 346 + col) <= 46018) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 46021 && (row * 346 + col) <= 46058) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46059 && (row * 346 + col) <= 46061) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46062 && (row * 346 + col) <= 46072) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46075 && (row * 346 + col) <= 46078) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46079 && (row * 346 + col) <= 46080) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46081 && (row * 346 + col) <= 46085) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46086 && (row * 346 + col) <= 46087) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46088 && (row * 346 + col) <= 46089) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46090 && (row * 346 + col) <= 46091) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46092 && (row * 346 + col) <= 46092) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46093 && (row * 346 + col) <= 46094) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46095 && (row * 346 + col) <= 46095) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46096 && (row * 346 + col) <= 46097) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46098 && (row * 346 + col) <= 46098) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46099 && (row * 346 + col) <= 46100) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46101 && (row * 346 + col) <= 46102) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46103 && (row * 346 + col) <= 46104) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46105 && (row * 346 + col) <= 46108) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46111 && (row * 346 + col) <= 46140) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46153 && (row * 346 + col) <= 46158) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46165 && (row * 346 + col) <= 46176) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46192 && (row * 346 + col) <= 46196) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46208 && (row * 346 + col) <= 46224) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46240 && (row * 346 + col) <= 46242) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46249 && (row * 346 + col) <= 46251) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46258 && (row * 346 + col) <= 46260) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46276 && (row * 346 + col) <= 46281) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46288 && (row * 346 + col) <= 46293) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46300 && (row * 346 + col) <= 46302) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46312 && (row * 346 + col) <= 46323) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46324 && (row * 346 + col) <= 46326) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46327 && (row * 346 + col) <= 46360) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46363 && (row * 346 + col) <= 46364) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 46367 && (row * 346 + col) <= 46404) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46405 && (row * 346 + col) <= 46407) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46408 && (row * 346 + col) <= 46418) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46421 && (row * 346 + col) <= 46425) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46426 && (row * 346 + col) <= 46428) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46429 && (row * 346 + col) <= 46431) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46432 && (row * 346 + col) <= 46433) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46434 && (row * 346 + col) <= 46435) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46436 && (row * 346 + col) <= 46440) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46441 && (row * 346 + col) <= 46441) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46442 && (row * 346 + col) <= 46445) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46446 && (row * 346 + col) <= 46448) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46449 && (row * 346 + col) <= 46450) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46451 && (row * 346 + col) <= 46454) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46457 && (row * 346 + col) <= 46486) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46499 && (row * 346 + col) <= 46504) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46511 && (row * 346 + col) <= 46522) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46538 && (row * 346 + col) <= 46543) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46553 && (row * 346 + col) <= 46570) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46586 && (row * 346 + col) <= 46588) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46595 && (row * 346 + col) <= 46597) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46604 && (row * 346 + col) <= 46606) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46622 && (row * 346 + col) <= 46627) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46634 && (row * 346 + col) <= 46639) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46646 && (row * 346 + col) <= 46648) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46658 && (row * 346 + col) <= 46669) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46670 && (row * 346 + col) <= 46672) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46673 && (row * 346 + col) <= 46706) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46709 && (row * 346 + col) <= 46710) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 46713 && (row * 346 + col) <= 46750) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46751 && (row * 346 + col) <= 46753) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46754 && (row * 346 + col) <= 46764) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46767 && (row * 346 + col) <= 46773) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46774 && (row * 346 + col) <= 46775) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46776 && (row * 346 + col) <= 46777) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46778 && (row * 346 + col) <= 46779) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46780 && (row * 346 + col) <= 46781) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46782 && (row * 346 + col) <= 46783) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46784 && (row * 346 + col) <= 46784) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46785 && (row * 346 + col) <= 46786) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46787 && (row * 346 + col) <= 46787) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46788 && (row * 346 + col) <= 46789) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46790 && (row * 346 + col) <= 46790) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46791 && (row * 346 + col) <= 46792) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46793 && (row * 346 + col) <= 46794) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46795 && (row * 346 + col) <= 46796) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46797 && (row * 346 + col) <= 46800) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 46803 && (row * 346 + col) <= 46832) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46845 && (row * 346 + col) <= 46850) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46857 && (row * 346 + col) <= 46868) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46884 && (row * 346 + col) <= 46889) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46899 && (row * 346 + col) <= 46916) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46932 && (row * 346 + col) <= 46934) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46941 && (row * 346 + col) <= 46943) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46950 && (row * 346 + col) <= 46952) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46968 && (row * 346 + col) <= 46973) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46980 && (row * 346 + col) <= 46985) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 46992 && (row * 346 + col) <= 46994) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47004 && (row * 346 + col) <= 47015) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47016 && (row * 346 + col) <= 47018) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47019 && (row * 346 + col) <= 47052) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47055 && (row * 346 + col) <= 47056) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 47059 && (row * 346 + col) <= 47096) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47097 && (row * 346 + col) <= 47099) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47100 && (row * 346 + col) <= 47110) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47113 && (row * 346 + col) <= 47119) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47120 && (row * 346 + col) <= 47121) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47122 && (row * 346 + col) <= 47123) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47124 && (row * 346 + col) <= 47125) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47126 && (row * 346 + col) <= 47127) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47128 && (row * 346 + col) <= 47129) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47130 && (row * 346 + col) <= 47130) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47131 && (row * 346 + col) <= 47132) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47133 && (row * 346 + col) <= 47133) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47134 && (row * 346 + col) <= 47135) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47136 && (row * 346 + col) <= 47136) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47137 && (row * 346 + col) <= 47138) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47139 && (row * 346 + col) <= 47140) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47141 && (row * 346 + col) <= 47142) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47143 && (row * 346 + col) <= 47146) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47149 && (row * 346 + col) <= 47178) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47185 && (row * 346 + col) <= 47196) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47203 && (row * 346 + col) <= 47214) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47221 && (row * 346 + col) <= 47223) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47230 && (row * 346 + col) <= 47237) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47243 && (row * 346 + col) <= 47262) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47269 && (row * 346 + col) <= 47271) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47278 && (row * 346 + col) <= 47280) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47287 && (row * 346 + col) <= 47289) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47296 && (row * 346 + col) <= 47298) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47305 && (row * 346 + col) <= 47307) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47314 && (row * 346 + col) <= 47319) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47326 && (row * 346 + col) <= 47331) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47338 && (row * 346 + col) <= 47343) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47350 && (row * 346 + col) <= 47361) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47362 && (row * 346 + col) <= 47364) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47365 && (row * 346 + col) <= 47398) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47401 && (row * 346 + col) <= 47402) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 47405 && (row * 346 + col) <= 47442) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47443 && (row * 346 + col) <= 47445) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47446 && (row * 346 + col) <= 47456) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47459 && (row * 346 + col) <= 47462) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47463 && (row * 346 + col) <= 47464) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47465 && (row * 346 + col) <= 47465) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47466 && (row * 346 + col) <= 47467) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47468 && (row * 346 + col) <= 47469) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47470 && (row * 346 + col) <= 47471) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47472 && (row * 346 + col) <= 47473) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47474 && (row * 346 + col) <= 47475) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47476 && (row * 346 + col) <= 47476) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47477 && (row * 346 + col) <= 47478) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47479 && (row * 346 + col) <= 47479) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47480 && (row * 346 + col) <= 47481) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47482 && (row * 346 + col) <= 47482) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47483 && (row * 346 + col) <= 47484) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47485 && (row * 346 + col) <= 47486) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47487 && (row * 346 + col) <= 47488) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47489 && (row * 346 + col) <= 47492) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47495 && (row * 346 + col) <= 47524) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47531 && (row * 346 + col) <= 47542) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47549 && (row * 346 + col) <= 47560) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47567 && (row * 346 + col) <= 47569) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47576 && (row * 346 + col) <= 47583) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47589 && (row * 346 + col) <= 47608) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47615 && (row * 346 + col) <= 47617) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47624 && (row * 346 + col) <= 47626) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47633 && (row * 346 + col) <= 47635) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47642 && (row * 346 + col) <= 47644) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47651 && (row * 346 + col) <= 47653) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47660 && (row * 346 + col) <= 47665) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47672 && (row * 346 + col) <= 47677) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47684 && (row * 346 + col) <= 47689) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47696 && (row * 346 + col) <= 47707) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47708 && (row * 346 + col) <= 47710) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47711 && (row * 346 + col) <= 47744) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47747 && (row * 346 + col) <= 47748) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 47751 && (row * 346 + col) <= 47788) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47789 && (row * 346 + col) <= 47791) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47792 && (row * 346 + col) <= 47802) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47805 && (row * 346 + col) <= 47808) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47809 && (row * 346 + col) <= 47813) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47814 && (row * 346 + col) <= 47815) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47816 && (row * 346 + col) <= 47817) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47818 && (row * 346 + col) <= 47819) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47820 && (row * 346 + col) <= 47821) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47822 && (row * 346 + col) <= 47822) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47823 && (row * 346 + col) <= 47824) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47825 && (row * 346 + col) <= 47825) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47826 && (row * 346 + col) <= 47827) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47828 && (row * 346 + col) <= 47828) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47829 && (row * 346 + col) <= 47830) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47831 && (row * 346 + col) <= 47832) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47833 && (row * 346 + col) <= 47834) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47835 && (row * 346 + col) <= 47838) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 47841 && (row * 346 + col) <= 47870) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47877 && (row * 346 + col) <= 47888) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47895 && (row * 346 + col) <= 47906) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47913 && (row * 346 + col) <= 47915) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47922 && (row * 346 + col) <= 47929) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47935 && (row * 346 + col) <= 47954) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47961 && (row * 346 + col) <= 47963) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47970 && (row * 346 + col) <= 47972) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47979 && (row * 346 + col) <= 47981) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47988 && (row * 346 + col) <= 47990) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 47997 && (row * 346 + col) <= 47999) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48006 && (row * 346 + col) <= 48011) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48018 && (row * 346 + col) <= 48023) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48030 && (row * 346 + col) <= 48035) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48042 && (row * 346 + col) <= 48053) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48054 && (row * 346 + col) <= 48056) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48057 && (row * 346 + col) <= 48090) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48093 && (row * 346 + col) <= 48094) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 48097 && (row * 346 + col) <= 48134) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48135 && (row * 346 + col) <= 48137) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48138 && (row * 346 + col) <= 48148) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48152 && (row * 346 + col) <= 48183) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48187 && (row * 346 + col) <= 48216) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48223 && (row * 346 + col) <= 48234) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48241 && (row * 346 + col) <= 48252) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48259 && (row * 346 + col) <= 48261) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48268 && (row * 346 + col) <= 48275) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48281 && (row * 346 + col) <= 48300) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48307 && (row * 346 + col) <= 48309) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48316 && (row * 346 + col) <= 48318) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48325 && (row * 346 + col) <= 48327) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48334 && (row * 346 + col) <= 48336) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48343 && (row * 346 + col) <= 48345) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48352 && (row * 346 + col) <= 48357) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48364 && (row * 346 + col) <= 48369) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48376 && (row * 346 + col) <= 48381) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48388 && (row * 346 + col) <= 48399) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48400 && (row * 346 + col) <= 48402) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48403 && (row * 346 + col) <= 48436) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48439 && (row * 346 + col) <= 48440) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 48443 && (row * 346 + col) <= 48480) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48481 && (row * 346 + col) <= 48483) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48484 && (row * 346 + col) <= 48495) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48498 && (row * 346 + col) <= 48529) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48532 && (row * 346 + col) <= 48562) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48569 && (row * 346 + col) <= 48580) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48587 && (row * 346 + col) <= 48598) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48605 && (row * 346 + col) <= 48607) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48614 && (row * 346 + col) <= 48621) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48627 && (row * 346 + col) <= 48646) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48653 && (row * 346 + col) <= 48655) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48662 && (row * 346 + col) <= 48664) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48671 && (row * 346 + col) <= 48673) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48680 && (row * 346 + col) <= 48682) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48689 && (row * 346 + col) <= 48691) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48698 && (row * 346 + col) <= 48703) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48710 && (row * 346 + col) <= 48715) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48722 && (row * 346 + col) <= 48727) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48734 && (row * 346 + col) <= 48745) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48746 && (row * 346 + col) <= 48748) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48749 && (row * 346 + col) <= 48782) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48785 && (row * 346 + col) <= 48786) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 48789 && (row * 346 + col) <= 48826) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48827 && (row * 346 + col) <= 48829) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48830 && (row * 346 + col) <= 48841) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48844 && (row * 346 + col) <= 48875) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 48878 && (row * 346 + col) <= 48908) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48915 && (row * 346 + col) <= 48926) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48933 && (row * 346 + col) <= 48944) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48951 && (row * 346 + col) <= 48953) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48960 && (row * 346 + col) <= 48967) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48973 && (row * 346 + col) <= 48992) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 48999 && (row * 346 + col) <= 49001) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49008 && (row * 346 + col) <= 49010) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49017 && (row * 346 + col) <= 49019) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49026 && (row * 346 + col) <= 49028) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49035 && (row * 346 + col) <= 49037) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49044 && (row * 346 + col) <= 49049) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49056 && (row * 346 + col) <= 49061) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49068 && (row * 346 + col) <= 49073) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49080 && (row * 346 + col) <= 49091) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49092 && (row * 346 + col) <= 49094) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49095 && (row * 346 + col) <= 49128) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49131 && (row * 346 + col) <= 49132) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 49135 && (row * 346 + col) <= 49172) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49173 && (row * 346 + col) <= 49175) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49176 && (row * 346 + col) <= 49187) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49191 && (row * 346 + col) <= 49220) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49224 && (row * 346 + col) <= 49237) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49242 && (row * 346 + col) <= 49254) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49261 && (row * 346 + col) <= 49272) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49279 && (row * 346 + col) <= 49290) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49297 && (row * 346 + col) <= 49299) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49306 && (row * 346 + col) <= 49313) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49319 && (row * 346 + col) <= 49338) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49345 && (row * 346 + col) <= 49347) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49354 && (row * 346 + col) <= 49356) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49363 && (row * 346 + col) <= 49365) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49372 && (row * 346 + col) <= 49374) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49381 && (row * 346 + col) <= 49383) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49390 && (row * 346 + col) <= 49395) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49402 && (row * 346 + col) <= 49407) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49414 && (row * 346 + col) <= 49419) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49426 && (row * 346 + col) <= 49437) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49438 && (row * 346 + col) <= 49440) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49441 && (row * 346 + col) <= 49474) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49477 && (row * 346 + col) <= 49478) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 49481 && (row * 346 + col) <= 49518) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49519 && (row * 346 + col) <= 49521) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49522 && (row * 346 + col) <= 49534) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49537 && (row * 346 + col) <= 49566) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49569 && (row * 346 + col) <= 49583) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49588 && (row * 346 + col) <= 49600) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49607 && (row * 346 + col) <= 49618) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49625 && (row * 346 + col) <= 49636) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49643 && (row * 346 + col) <= 49645) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49652 && (row * 346 + col) <= 49659) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49665 && (row * 346 + col) <= 49684) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49691 && (row * 346 + col) <= 49693) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49700 && (row * 346 + col) <= 49702) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49709 && (row * 346 + col) <= 49711) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49718 && (row * 346 + col) <= 49720) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49727 && (row * 346 + col) <= 49729) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49736 && (row * 346 + col) <= 49741) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49748 && (row * 346 + col) <= 49753) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49760 && (row * 346 + col) <= 49765) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49772 && (row * 346 + col) <= 49783) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49784 && (row * 346 + col) <= 49786) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49787 && (row * 346 + col) <= 49820) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49823 && (row * 346 + col) <= 49824) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 49827 && (row * 346 + col) <= 49864) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49865 && (row * 346 + col) <= 49867) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49868 && (row * 346 + col) <= 49880) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49884 && (row * 346 + col) <= 49911) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 49915 && (row * 346 + col) <= 49929) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49934 && (row * 346 + col) <= 49946) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49953 && (row * 346 + col) <= 49964) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49971 && (row * 346 + col) <= 49982) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49989 && (row * 346 + col) <= 49991) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 49998 && (row * 346 + col) <= 50005) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50011 && (row * 346 + col) <= 50030) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50037 && (row * 346 + col) <= 50039) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50046 && (row * 346 + col) <= 50048) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50055 && (row * 346 + col) <= 50057) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50064 && (row * 346 + col) <= 50066) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50073 && (row * 346 + col) <= 50075) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50082 && (row * 346 + col) <= 50087) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50094 && (row * 346 + col) <= 50099) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50106 && (row * 346 + col) <= 50111) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50118 && (row * 346 + col) <= 50129) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50130 && (row * 346 + col) <= 50132) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50133 && (row * 346 + col) <= 50166) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50169 && (row * 346 + col) <= 50170) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 50173 && (row * 346 + col) <= 50210) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50211 && (row * 346 + col) <= 50213) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50214 && (row * 346 + col) <= 50227) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50231 && (row * 346 + col) <= 50256) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50260 && (row * 346 + col) <= 50275) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50280 && (row * 346 + col) <= 50292) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50299 && (row * 346 + col) <= 50310) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50326 && (row * 346 + col) <= 50328) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50335 && (row * 346 + col) <= 50337) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50344 && (row * 346 + col) <= 50351) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50357 && (row * 346 + col) <= 50376) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50383 && (row * 346 + col) <= 50385) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50392 && (row * 346 + col) <= 50394) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50410 && (row * 346 + col) <= 50412) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50419 && (row * 346 + col) <= 50421) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50428 && (row * 346 + col) <= 50430) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50443 && (row * 346 + col) <= 50445) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50452 && (row * 346 + col) <= 50457) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50464 && (row * 346 + col) <= 50475) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50476 && (row * 346 + col) <= 50478) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50479 && (row * 346 + col) <= 50512) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50515 && (row * 346 + col) <= 50516) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 50519 && (row * 346 + col) <= 50556) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50557 && (row * 346 + col) <= 50559) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50560 && (row * 346 + col) <= 50574) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50578 && (row * 346 + col) <= 50601) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50605 && (row * 346 + col) <= 50638) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50645 && (row * 346 + col) <= 50656) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50672 && (row * 346 + col) <= 50674) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50681 && (row * 346 + col) <= 50683) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50690 && (row * 346 + col) <= 50697) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50703 && (row * 346 + col) <= 50722) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50729 && (row * 346 + col) <= 50731) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50738 && (row * 346 + col) <= 50740) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50756 && (row * 346 + col) <= 50758) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50765 && (row * 346 + col) <= 50767) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50774 && (row * 346 + col) <= 50776) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50789 && (row * 346 + col) <= 50791) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50798 && (row * 346 + col) <= 50803) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50810 && (row * 346 + col) <= 50821) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50822 && (row * 346 + col) <= 50824) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50825 && (row * 346 + col) <= 50858) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50861 && (row * 346 + col) <= 50862) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 50865 && (row * 346 + col) <= 50902) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50903 && (row * 346 + col) <= 50905) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50906 && (row * 346 + col) <= 50921) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50925 && (row * 346 + col) <= 50946) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 50950 && (row * 346 + col) <= 50984) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 50991 && (row * 346 + col) <= 51002) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51018 && (row * 346 + col) <= 51020) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51027 && (row * 346 + col) <= 51029) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51036 && (row * 346 + col) <= 51043) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51049 && (row * 346 + col) <= 51068) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51075 && (row * 346 + col) <= 51077) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51084 && (row * 346 + col) <= 51086) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51102 && (row * 346 + col) <= 51104) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51111 && (row * 346 + col) <= 51113) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51120 && (row * 346 + col) <= 51122) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51135 && (row * 346 + col) <= 51137) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51144 && (row * 346 + col) <= 51149) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51156 && (row * 346 + col) <= 51167) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51168 && (row * 346 + col) <= 51170) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51171 && (row * 346 + col) <= 51204) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51207 && (row * 346 + col) <= 51208) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 51211 && (row * 346 + col) <= 51248) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51249 && (row * 346 + col) <= 51251) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51252 && (row * 346 + col) <= 51268) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51272 && (row * 346 + col) <= 51291) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51295 && (row * 346 + col) <= 51513) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51514 && (row * 346 + col) <= 51516) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51517 && (row * 346 + col) <= 51550) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51553 && (row * 346 + col) <= 51554) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 51557 && (row * 346 + col) <= 51594) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51595 && (row * 346 + col) <= 51597) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51598 && (row * 346 + col) <= 51615) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51619 && (row * 346 + col) <= 51636) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51640 && (row * 346 + col) <= 51859) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51860 && (row * 346 + col) <= 51862) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51863 && (row * 346 + col) <= 51896) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51899 && (row * 346 + col) <= 51900) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 51903 && (row * 346 + col) <= 51940) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51941 && (row * 346 + col) <= 51943) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51944 && (row * 346 + col) <= 51962) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 51967 && (row * 346 + col) <= 51980) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 51985 && (row * 346 + col) <= 52205) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52206 && (row * 346 + col) <= 52208) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 52209 && (row * 346 + col) <= 52242) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52245 && (row * 346 + col) <= 52246) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 52249 && (row * 346 + col) <= 52286) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52287 && (row * 346 + col) <= 52289) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 52290 && (row * 346 + col) <= 52309) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52316 && (row * 346 + col) <= 52323) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 52330 && (row * 346 + col) <= 52551) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52552 && (row * 346 + col) <= 52554) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 52555 && (row * 346 + col) <= 52588) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52591 && (row * 346 + col) <= 52592) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 52595 && (row * 346 + col) <= 52632) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52633 && (row * 346 + col) <= 52635) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 52636 && (row * 346 + col) <= 52657) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52674 && (row * 346 + col) <= 52897) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52898 && (row * 346 + col) <= 52900) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 52901 && (row * 346 + col) <= 52934) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52937 && (row * 346 + col) <= 52938) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 52941 && (row * 346 + col) <= 52978) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 52979 && (row * 346 + col) <= 52981) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 52982 && (row * 346 + col) <= 53006) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53017 && (row * 346 + col) <= 53243) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53244 && (row * 346 + col) <= 53246) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 53247 && (row * 346 + col) <= 53280) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53283 && (row * 346 + col) <= 53284) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 53287 && (row * 346 + col) <= 53324) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53325 && (row * 346 + col) <= 53327) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 53328 && (row * 346 + col) <= 53589) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53590 && (row * 346 + col) <= 53592) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 53593 && (row * 346 + col) <= 53626) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53629 && (row * 346 + col) <= 53630) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 53633 && (row * 346 + col) <= 53670) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53671 && (row * 346 + col) <= 53673) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 53674 && (row * 346 + col) <= 53935) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53936 && (row * 346 + col) <= 53938) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 53939 && (row * 346 + col) <= 53972) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 53975 && (row * 346 + col) <= 53976) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 53979 && (row * 346 + col) <= 54016) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54017 && (row * 346 + col) <= 54019) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 54020 && (row * 346 + col) <= 54281) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54282 && (row * 346 + col) <= 54284) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 54285 && (row * 346 + col) <= 54318) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54321 && (row * 346 + col) <= 54322) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 54325 && (row * 346 + col) <= 54362) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54363 && (row * 346 + col) <= 54365) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 54366 && (row * 346 + col) <= 54627) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54628 && (row * 346 + col) <= 54630) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 54631 && (row * 346 + col) <= 54664) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54667 && (row * 346 + col) <= 54668) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 54671 && (row * 346 + col) <= 54708) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54709 && (row * 346 + col) <= 54711) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 54712 && (row * 346 + col) <= 54973) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 54974 && (row * 346 + col) <= 54976) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 54977 && (row * 346 + col) <= 55010) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55013 && (row * 346 + col) <= 55014) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 55017 && (row * 346 + col) <= 55054) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55055 && (row * 346 + col) <= 55057) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 55058 && (row * 346 + col) <= 55319) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55320 && (row * 346 + col) <= 55322) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 55323 && (row * 346 + col) <= 55356) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55359 && (row * 346 + col) <= 55360) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 55363 && (row * 346 + col) <= 55400) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55401 && (row * 346 + col) <= 55403) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 55404 && (row * 346 + col) <= 55665) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55666 && (row * 346 + col) <= 55668) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 55669 && (row * 346 + col) <= 55702) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55705 && (row * 346 + col) <= 55706) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 55709 && (row * 346 + col) <= 55746) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 55747 && (row * 346 + col) <= 55749) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 55750 && (row * 346 + col) <= 56011) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56012 && (row * 346 + col) <= 56014) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 56015 && (row * 346 + col) <= 56048) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56051 && (row * 346 + col) <= 56052) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 56055 && (row * 346 + col) <= 56092) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56093 && (row * 346 + col) <= 56095) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 56096 && (row * 346 + col) <= 56357) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56358 && (row * 346 + col) <= 56360) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 56361 && (row * 346 + col) <= 56394) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56397 && (row * 346 + col) <= 56398) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 56401 && (row * 346 + col) <= 56438) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56439 && (row * 346 + col) <= 56441) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 56442 && (row * 346 + col) <= 56703) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56704 && (row * 346 + col) <= 56706) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 56707 && (row * 346 + col) <= 56740) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56743 && (row * 346 + col) <= 56744) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 56747 && (row * 346 + col) <= 56784) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 56785 && (row * 346 + col) <= 56787) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 56788 && (row * 346 + col) <= 57049) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 57050 && (row * 346 + col) <= 57052) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 57053 && (row * 346 + col) <= 57086) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 57089 && (row * 346 + col) <= 57090) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 57093 && (row * 346 + col) <= 57130) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 57131 && (row * 346 + col) <= 57398) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 57399 && (row * 346 + col) <= 57432) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 57435 && (row * 346 + col) <= 57436) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 57443 && (row * 346 + col) <= 57476) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 57477 && (row * 346 + col) <= 57744) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 57745 && (row * 346 + col) <= 57774) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 57781 && (row * 346 + col) <= 57782) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 57789 && (row * 346 + col) <= 57822) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 57823 && (row * 346 + col) <= 58090) color_data <= 12'b110011001100; else
        if ((row * 346 + col) >= 58091 && (row * 346 + col) <= 58120) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 58127 && (row * 346 + col) <= 58132) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 58135 && (row * 346 + col) <= 58466) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 58469 && (row * 346 + col) <= 58478) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 58481 && (row * 346 + col) <= 58812) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 58815 && (row * 346 + col) <= 58824) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 58827 && (row * 346 + col) <= 59158) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 59161 && (row * 346 + col) <= 59170) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 59173 && (row * 346 + col) <= 59504) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 59507 && (row * 346 + col) <= 59516) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 59519 && (row * 346 + col) <= 59850) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 59853 && (row * 346 + col) <= 59862) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 59865 && (row * 346 + col) <= 60196) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 60199 && (row * 346 + col) <= 60208) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 60215 && (row * 346 + col) <= 60538) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 60545 && (row * 346 + col) <= 60554) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 60561 && (row * 346 + col) <= 60884) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 60891 && (row * 346 + col) <= 60904) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 60907 && (row * 346 + col) <= 61230) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 61233 && (row * 346 + col) <= 61250) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 61253 && (row * 346 + col) <= 61576) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 61579 && (row * 346 + col) <= 61596) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 61607 && (row * 346 + col) <= 61914) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 61925 && (row * 346 + col) <= 61942) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 61953 && (row * 346 + col) <= 62260) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 62271 && (row * 346 + col) <= 62296) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 62299 && (row * 346 + col) <= 62606) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 62609 && (row * 346 + col) <= 62642) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 62645 && (row * 346 + col) <= 62952) color_data <= 12'b101010101010; else
        if ((row * 346 + col) >= 62955 && (row * 346 + col) <= 62988) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 63301 && (row * 346 + col) <= 63334) color_data <= 12'b111111111111; else
        if ((row * 346 + col) >= 63647 && (row * 346 + col) < 64010) color_data <= 12'b111111111111; else
        color_data <= 12'b000000000000;
    end
endmodule