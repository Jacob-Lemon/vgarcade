`timescale 1ns / 1ps
module background_rom (
    input wire clk,
    input wire [8:0] row,
    input wire [9:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ( {row,col} >= 000000 && {row,col} <= 000131) color_data <= 12'b111111110000; else
        if ( {row,col} >= 000132 && {row,col} <= 000639) color_data <= 12'b000010101110; else
        if ( {row,col} >= 000640 && {row,col} <= 000771) color_data <= 12'b111111110000; else
        if ( {row,col} >= 000772 && {row,col} <= 001279) color_data <= 12'b000010101110; else
        if ( {row,col} >= 001280 && {row,col} <= 001411) color_data <= 12'b111111110000; else
        if ( {row,col} >= 001412 && {row,col} <= 001919) color_data <= 12'b000010101110; else
        if ( {row,col} >= 001920 && {row,col} <= 002051) color_data <= 12'b111111110000; else
        if ( {row,col} >= 002052 && {row,col} <= 002559) color_data <= 12'b000010101110; else
        if ( {row,col} >= 002560 && {row,col} <= 002691) color_data <= 12'b111111110000; else
        if ( {row,col} >= 002692 && {row,col} <= 003199) color_data <= 12'b000010101110; else
        if ( {row,col} >= 003200 && {row,col} <= 003331) color_data <= 12'b111111110000; else
        if ( {row,col} >= 003332 && {row,col} <= 003839) color_data <= 12'b000010101110; else
        if ( {row,col} >= 003840 && {row,col} <= 003971) color_data <= 12'b111111110000; else
        if ( {row,col} >= 003972 && {row,col} <= 004479) color_data <= 12'b000010101110; else
        if ( {row,col} >= 004480 && {row,col} <= 004611) color_data <= 12'b111111110000; else
        if ( {row,col} >= 004612 && {row,col} <= 005119) color_data <= 12'b000010101110; else
        if ( {row,col} >= 005120 && {row,col} <= 005251) color_data <= 12'b111111110000; else
        if ( {row,col} >= 005252 && {row,col} <= 005759) color_data <= 12'b000010101110; else
        if ( {row,col} >= 005760 && {row,col} <= 005890) color_data <= 12'b111111110000; else
        if ( {row,col} >= 005891 && {row,col} <= 006399) color_data <= 12'b000010101110; else
        if ( {row,col} >= 006400 && {row,col} <= 006530) color_data <= 12'b111111110000; else
        if ( {row,col} >= 006531 && {row,col} <= 007039) color_data <= 12'b000010101110; else
        if ( {row,col} >= 007040 && {row,col} <= 007170) color_data <= 12'b111111110000; else
        if ( {row,col} >= 007171 && {row,col} <= 007679) color_data <= 12'b000010101110; else
        if ( {row,col} >= 007680 && {row,col} <= 007810) color_data <= 12'b111111110000; else
        if ( {row,col} >= 007811 && {row,col} <= 008319) color_data <= 12'b000010101110; else
        if ( {row,col} >= 008320 && {row,col} <= 008450) color_data <= 12'b111111110000; else
        if ( {row,col} >= 008451 && {row,col} <= 008959) color_data <= 12'b000010101110; else
        if ( {row,col} >= 008960 && {row,col} <= 009090) color_data <= 12'b111111110000; else
        if ( {row,col} >= 009091 && {row,col} <= 009507) color_data <= 12'b000010101110; else
        if ( {row,col} >= 009508 && {row,col} <= 009514) color_data <= 12'b111111111111; else
        if ( {row,col} >= 009515 && {row,col} <= 009525) color_data <= 12'b000010101110; else
        if ( {row,col} >= 009526 && {row,col} <= 009533) color_data <= 12'b111111111111; else
        if ( {row,col} >= 009534 && {row,col} <= 009599) color_data <= 12'b000010101110; else
        if ( {row,col} >= 009600 && {row,col} <= 009730) color_data <= 12'b111111110000; else
        if ( {row,col} >= 009731 && {row,col} <= 010143) color_data <= 12'b000010101110; else
        if ( {row,col} >= 010144 && {row,col} <= 010157) color_data <= 12'b111111111111; else
        if ( {row,col} >= 010158 && {row,col} <= 010162) color_data <= 12'b000010101110; else
        if ( {row,col} >= 010163 && {row,col} <= 010177) color_data <= 12'b111111111111; else
        if ( {row,col} >= 010178 && {row,col} <= 010239) color_data <= 12'b000010101110; else
        if ( {row,col} >= 010240 && {row,col} <= 010370) color_data <= 12'b111111110000; else
        if ( {row,col} >= 010371 && {row,col} <= 010765) color_data <= 12'b000010101110; else
        if ( {row,col} >= 010766 && {row,col} <= 010776) color_data <= 12'b111111111111; else
        if ( {row,col} >= 010777 && {row,col} <= 010781) color_data <= 12'b000010101110; else
        if ( {row,col} >= 010782 && {row,col} <= 010819) color_data <= 12'b111111111111; else
        if ( {row,col} >= 010820 && {row,col} <= 010879) color_data <= 12'b000010101110; else
        if ( {row,col} >= 010880 && {row,col} <= 011010) color_data <= 12'b111111110000; else
        if ( {row,col} >= 011011 && {row,col} <= 011402) color_data <= 12'b000010101110; else
        if ( {row,col} >= 011403 && {row,col} <= 011461) color_data <= 12'b111111111111; else
        if ( {row,col} >= 011462 && {row,col} <= 011519) color_data <= 12'b000010101110; else
        if ( {row,col} >= 011520 && {row,col} <= 011649) color_data <= 12'b111111110000; else
        if ( {row,col} >= 011650 && {row,col} <= 012040) color_data <= 12'b000010101110; else
        if ( {row,col} >= 012041 && {row,col} <= 012102) color_data <= 12'b111111111111; else
        if ( {row,col} >= 012103 && {row,col} <= 012159) color_data <= 12'b000010101110; else
        if ( {row,col} >= 012160 && {row,col} <= 012289) color_data <= 12'b111111110000; else
        if ( {row,col} >= 012290 && {row,col} <= 012662) color_data <= 12'b000010101110; else
        if ( {row,col} >= 012663 && {row,col} <= 012676) color_data <= 12'b111111111111; else
        if ( {row,col} >= 012677 && {row,col} <= 012678) color_data <= 12'b000010101110; else
        if ( {row,col} >= 012679 && {row,col} <= 012743) color_data <= 12'b111111111111; else
        if ( {row,col} >= 012744 && {row,col} <= 012799) color_data <= 12'b000010101110; else
        if ( {row,col} >= 012800 && {row,col} <= 012929) color_data <= 12'b111111110000; else
        if ( {row,col} >= 012930 && {row,col} <= 013299) color_data <= 12'b000010101110; else
        if ( {row,col} >= 013300 && {row,col} <= 013384) color_data <= 12'b111111111111; else
        if ( {row,col} >= 013385 && {row,col} <= 013439) color_data <= 12'b000010101110; else
        if ( {row,col} >= 013440 && {row,col} <= 013569) color_data <= 12'b111111110000; else
        if ( {row,col} >= 013570 && {row,col} <= 013937) color_data <= 12'b000010101110; else
        if ( {row,col} >= 013938 && {row,col} <= 014026) color_data <= 12'b111111111111; else
        if ( {row,col} >= 014027 && {row,col} <= 014079) color_data <= 12'b000010101110; else
        if ( {row,col} >= 014080 && {row,col} <= 014209) color_data <= 12'b111111110000; else
        if ( {row,col} >= 014210 && {row,col} <= 014575) color_data <= 12'b000010101110; else
        if ( {row,col} >= 014576 && {row,col} <= 014668) color_data <= 12'b111111111111; else
        if ( {row,col} >= 014669 && {row,col} <= 014719) color_data <= 12'b000010101110; else
        if ( {row,col} >= 014720 && {row,col} <= 014849) color_data <= 12'b111111110000; else
        if ( {row,col} >= 014850 && {row,col} <= 015214) color_data <= 12'b000010101110; else
        if ( {row,col} >= 015215 && {row,col} <= 015310) color_data <= 12'b111111111111; else
        if ( {row,col} >= 015311 && {row,col} <= 015359) color_data <= 12'b000010101110; else
        if ( {row,col} >= 015360 && {row,col} <= 015488) color_data <= 12'b111111110000; else
        if ( {row,col} >= 015489 && {row,col} <= 015853) color_data <= 12'b000010101110; else
        if ( {row,col} >= 015854 && {row,col} <= 015951) color_data <= 12'b111111111111; else
        if ( {row,col} >= 015952 && {row,col} <= 015999) color_data <= 12'b000010101110; else
        if ( {row,col} >= 016000 && {row,col} <= 016128) color_data <= 12'b111111110000; else
        if ( {row,col} >= 016129 && {row,col} <= 016492) color_data <= 12'b000010101110; else
        if ( {row,col} >= 016493 && {row,col} <= 016592) color_data <= 12'b111111111111; else
        if ( {row,col} >= 016593 && {row,col} <= 016639) color_data <= 12'b000010101110; else
        if ( {row,col} >= 016640 && {row,col} <= 016768) color_data <= 12'b111111110000; else
        if ( {row,col} >= 016769 && {row,col} <= 017131) color_data <= 12'b000010101110; else
        if ( {row,col} >= 017132 && {row,col} <= 017233) color_data <= 12'b111111111111; else
        if ( {row,col} >= 017234 && {row,col} <= 017279) color_data <= 12'b000010101110; else
        if ( {row,col} >= 017280 && {row,col} <= 017408) color_data <= 12'b111111110000; else
        if ( {row,col} >= 017409 && {row,col} <= 017771) color_data <= 12'b000010101110; else
        if ( {row,col} >= 017772 && {row,col} <= 017874) color_data <= 12'b111111111111; else
        if ( {row,col} >= 017875 && {row,col} <= 017919) color_data <= 12'b000010101110; else
        if ( {row,col} >= 017920 && {row,col} <= 018047) color_data <= 12'b111111110000; else
        if ( {row,col} >= 018048 && {row,col} <= 018410) color_data <= 12'b000010101110; else
        if ( {row,col} >= 018411 && {row,col} <= 018514) color_data <= 12'b111111111111; else
        if ( {row,col} >= 018515 && {row,col} <= 018559) color_data <= 12'b000010101110; else
        if ( {row,col} >= 018560 && {row,col} <= 018687) color_data <= 12'b111111110000; else
        if ( {row,col} >= 018688 && {row,col} <= 019050) color_data <= 12'b000010101110; else
        if ( {row,col} >= 019051 && {row,col} <= 019154) color_data <= 12'b111111111111; else
        if ( {row,col} >= 019155 && {row,col} <= 019199) color_data <= 12'b000010101110; else
        if ( {row,col} >= 019200 && {row,col} <= 019327) color_data <= 12'b111111110000; else
        if ( {row,col} >= 019328 && {row,col} <= 019690) color_data <= 12'b000010101110; else
        if ( {row,col} >= 019691 && {row,col} <= 019795) color_data <= 12'b111111111111; else
        if ( {row,col} >= 019796 && {row,col} <= 019839) color_data <= 12'b000010101110; else
        if ( {row,col} >= 019840 && {row,col} <= 019967) color_data <= 12'b111111110000; else
        if ( {row,col} >= 019968 && {row,col} <= 020326) color_data <= 12'b000010101110; else
        if ( {row,col} >= 020327 && {row,col} <= 020435) color_data <= 12'b111111111111; else
        if ( {row,col} >= 020436 && {row,col} <= 020479) color_data <= 12'b000010101110; else
        if ( {row,col} >= 020480 && {row,col} <= 020606) color_data <= 12'b111111110000; else
        if ( {row,col} >= 020607 && {row,col} <= 020964) color_data <= 12'b000010101110; else
        if ( {row,col} >= 020965 && {row,col} <= 021074) color_data <= 12'b111111111111; else
        if ( {row,col} >= 021075 && {row,col} <= 021119) color_data <= 12'b000010101110; else
        if ( {row,col} >= 021120 && {row,col} <= 021246) color_data <= 12'b111111110000; else
        if ( {row,col} >= 021247 && {row,col} <= 021602) color_data <= 12'b000010101110; else
        if ( {row,col} >= 021603 && {row,col} <= 021714) color_data <= 12'b111111111111; else
        if ( {row,col} >= 021715 && {row,col} <= 021759) color_data <= 12'b000010101110; else
        if ( {row,col} >= 021760 && {row,col} <= 021886) color_data <= 12'b111111110000; else
        if ( {row,col} >= 021887 && {row,col} <= 022240) color_data <= 12'b000010101110; else
        if ( {row,col} >= 022241 && {row,col} <= 022355) color_data <= 12'b111111111111; else
        if ( {row,col} >= 022356 && {row,col} <= 022399) color_data <= 12'b000010101110; else
        if ( {row,col} >= 022400 && {row,col} <= 022525) color_data <= 12'b111111110000; else
        if ( {row,col} >= 022526 && {row,col} <= 022880) color_data <= 12'b000010101110; else
        if ( {row,col} >= 022881 && {row,col} <= 022995) color_data <= 12'b111111111111; else
        if ( {row,col} >= 022996 && {row,col} <= 023039) color_data <= 12'b000010101110; else
        if ( {row,col} >= 023040 && {row,col} <= 023165) color_data <= 12'b111111110000; else
        if ( {row,col} >= 023166 && {row,col} <= 023519) color_data <= 12'b000010101110; else
        if ( {row,col} >= 023520 && {row,col} <= 023636) color_data <= 12'b111111111111; else
        if ( {row,col} >= 023637 && {row,col} <= 023679) color_data <= 12'b000010101110; else
        if ( {row,col} >= 023680 && {row,col} <= 023805) color_data <= 12'b111111110000; else
        if ( {row,col} >= 023806 && {row,col} <= 024158) color_data <= 12'b000010101110; else
        if ( {row,col} >= 024159 && {row,col} <= 024276) color_data <= 12'b111111111111; else
        if ( {row,col} >= 024277 && {row,col} <= 024319) color_data <= 12'b000010101110; else
        if ( {row,col} >= 024320 && {row,col} <= 024444) color_data <= 12'b111111110000; else
        if ( {row,col} >= 024445 && {row,col} <= 024798) color_data <= 12'b000010101110; else
        if ( {row,col} >= 024799 && {row,col} <= 024917) color_data <= 12'b111111111111; else
        if ( {row,col} >= 024918 && {row,col} <= 024959) color_data <= 12'b000010101110; else
        if ( {row,col} >= 024960 && {row,col} <= 025084) color_data <= 12'b111111110000; else
        if ( {row,col} >= 025085 && {row,col} <= 025438) color_data <= 12'b000010101110; else
        if ( {row,col} >= 025439 && {row,col} <= 025557) color_data <= 12'b111111111111; else
        if ( {row,col} >= 025558 && {row,col} <= 025599) color_data <= 12'b000010101110; else
        if ( {row,col} >= 025600 && {row,col} <= 025724) color_data <= 12'b111111110000; else
        if ( {row,col} >= 025725 && {row,col} <= 026078) color_data <= 12'b000010101110; else
        if ( {row,col} >= 026079 && {row,col} <= 026197) color_data <= 12'b111111111111; else
        if ( {row,col} >= 026198 && {row,col} <= 026239) color_data <= 12'b000010101110; else
        if ( {row,col} >= 026240 && {row,col} <= 026363) color_data <= 12'b111111110000; else
        if ( {row,col} >= 026364 && {row,col} <= 026718) color_data <= 12'b000010101110; else
        if ( {row,col} >= 026719 && {row,col} <= 026837) color_data <= 12'b111111111111; else
        if ( {row,col} >= 026838 && {row,col} <= 026879) color_data <= 12'b000010101110; else
        if ( {row,col} >= 026880 && {row,col} <= 027003) color_data <= 12'b111111110000; else
        if ( {row,col} >= 027004 && {row,col} <= 027359) color_data <= 12'b000010101110; else
        if ( {row,col} >= 027360 && {row,col} <= 027477) color_data <= 12'b111111111111; else
        if ( {row,col} >= 027478 && {row,col} <= 027519) color_data <= 12'b000010101110; else
        if ( {row,col} >= 027520 && {row,col} <= 027642) color_data <= 12'b111111110000; else
        if ( {row,col} >= 027643 && {row,col} <= 027999) color_data <= 12'b000010101110; else
        if ( {row,col} >= 028000 && {row,col} <= 028116) color_data <= 12'b111111111111; else
        if ( {row,col} >= 028117 && {row,col} <= 028159) color_data <= 12'b000010101110; else
        if ( {row,col} >= 028160 && {row,col} <= 028282) color_data <= 12'b111111110000; else
        if ( {row,col} >= 028283 && {row,col} <= 028640) color_data <= 12'b000010101110; else
        if ( {row,col} >= 028641 && {row,col} <= 028756) color_data <= 12'b111111111111; else
        if ( {row,col} >= 028757 && {row,col} <= 028799) color_data <= 12'b000010101110; else
        if ( {row,col} >= 028800 && {row,col} <= 028922) color_data <= 12'b111111110000; else
        if ( {row,col} >= 028923 && {row,col} <= 029281) color_data <= 12'b000010101110; else
        if ( {row,col} >= 029282 && {row,col} <= 029395) color_data <= 12'b111111111111; else
        if ( {row,col} >= 029396 && {row,col} <= 029439) color_data <= 12'b000010101110; else
        if ( {row,col} >= 029440 && {row,col} <= 029561) color_data <= 12'b111111110000; else
        if ( {row,col} >= 029562 && {row,col} <= 029923) color_data <= 12'b000010101110; else
        if ( {row,col} >= 029924 && {row,col} <= 030035) color_data <= 12'b111111111111; else
        if ( {row,col} >= 030036 && {row,col} <= 030079) color_data <= 12'b000010101110; else
        if ( {row,col} >= 030080 && {row,col} <= 030201) color_data <= 12'b111111110000; else
        if ( {row,col} >= 030202 && {row,col} <= 030562) color_data <= 12'b000010101110; else
        if ( {row,col} >= 030563 && {row,col} <= 030674) color_data <= 12'b111111111111; else
        if ( {row,col} >= 030675 && {row,col} <= 030719) color_data <= 12'b000010101110; else
        if ( {row,col} >= 030720 && {row,col} <= 030840) color_data <= 12'b111111110000; else
        if ( {row,col} >= 030841 && {row,col} <= 031202) color_data <= 12'b000010101110; else
        if ( {row,col} >= 031203 && {row,col} <= 031312) color_data <= 12'b111111111111; else
        if ( {row,col} >= 031313 && {row,col} <= 031359) color_data <= 12'b000010101110; else
        if ( {row,col} >= 031360 && {row,col} <= 031480) color_data <= 12'b111111110000; else
        if ( {row,col} >= 031481 && {row,col} <= 031842) color_data <= 12'b000010101110; else
        if ( {row,col} >= 031843 && {row,col} <= 031951) color_data <= 12'b111111111111; else
        if ( {row,col} >= 031952 && {row,col} <= 031999) color_data <= 12'b000010101110; else
        if ( {row,col} >= 032000 && {row,col} <= 032119) color_data <= 12'b111111110000; else
        if ( {row,col} >= 032120 && {row,col} <= 032482) color_data <= 12'b000010101110; else
        if ( {row,col} >= 032483 && {row,col} <= 032589) color_data <= 12'b111111111111; else
        if ( {row,col} >= 032590 && {row,col} <= 032639) color_data <= 12'b000010101110; else
        if ( {row,col} >= 032640 && {row,col} <= 032759) color_data <= 12'b111111110000; else
        if ( {row,col} >= 032760 && {row,col} <= 033122) color_data <= 12'b000010101110; else
        if ( {row,col} >= 033123 && {row,col} <= 033226) color_data <= 12'b111111111111; else
        if ( {row,col} >= 033227 && {row,col} <= 033279) color_data <= 12'b000010101110; else
        if ( {row,col} >= 033280 && {row,col} <= 033398) color_data <= 12'b111111110000; else
        if ( {row,col} >= 033399 && {row,col} <= 033762) color_data <= 12'b000010101110; else
        if ( {row,col} >= 033763 && {row,col} <= 033862) color_data <= 12'b111111111111; else
        if ( {row,col} >= 033863 && {row,col} <= 033919) color_data <= 12'b000010101110; else
        if ( {row,col} >= 033920 && {row,col} <= 034038) color_data <= 12'b111111110000; else
        if ( {row,col} >= 034039 && {row,col} <= 034402) color_data <= 12'b000010101110; else
        if ( {row,col} >= 034403 && {row,col} <= 034501) color_data <= 12'b111111111111; else
        if ( {row,col} >= 034502 && {row,col} <= 034559) color_data <= 12'b000010101110; else
        if ( {row,col} >= 034560 && {row,col} <= 034677) color_data <= 12'b111111110000; else
        if ( {row,col} >= 034678 && {row,col} <= 035043) color_data <= 12'b000010101110; else
        if ( {row,col} >= 035044 && {row,col} <= 035141) color_data <= 12'b111111111111; else
        if ( {row,col} >= 035142 && {row,col} <= 035199) color_data <= 12'b000010101110; else
        if ( {row,col} >= 035200 && {row,col} <= 035317) color_data <= 12'b111111110000; else
        if ( {row,col} >= 035318 && {row,col} <= 035684) color_data <= 12'b000010101110; else
        if ( {row,col} >= 035685 && {row,col} <= 035780) color_data <= 12'b111111111111; else
        if ( {row,col} >= 035781 && {row,col} <= 035839) color_data <= 12'b000010101110; else
        if ( {row,col} >= 035840 && {row,col} <= 035956) color_data <= 12'b111111110000; else
        if ( {row,col} >= 035957 && {row,col} <= 036325) color_data <= 12'b000010101110; else
        if ( {row,col} >= 036326 && {row,col} <= 036419) color_data <= 12'b111111111111; else
        if ( {row,col} >= 036420 && {row,col} <= 036479) color_data <= 12'b000010101110; else
        if ( {row,col} >= 036480 && {row,col} <= 036596) color_data <= 12'b111111110000; else
        if ( {row,col} >= 036597 && {row,col} <= 036967) color_data <= 12'b000010101110; else
        if ( {row,col} >= 036968 && {row,col} <= 037058) color_data <= 12'b111111111111; else
        if ( {row,col} >= 037059 && {row,col} <= 037119) color_data <= 12'b000010101110; else
        if ( {row,col} >= 037120 && {row,col} <= 037235) color_data <= 12'b111111110000; else
        if ( {row,col} >= 037236 && {row,col} <= 037609) color_data <= 12'b000010101110; else
        if ( {row,col} >= 037610 && {row,col} <= 037697) color_data <= 12'b111111111111; else
        if ( {row,col} >= 037698 && {row,col} <= 037759) color_data <= 12'b000010101110; else
        if ( {row,col} >= 037760 && {row,col} <= 037874) color_data <= 12'b111111110000; else
        if ( {row,col} >= 037875 && {row,col} <= 038253) color_data <= 12'b000010101110; else
        if ( {row,col} >= 038254 && {row,col} <= 038335) color_data <= 12'b111111111111; else
        if ( {row,col} >= 038336 && {row,col} <= 038399) color_data <= 12'b000010101110; else
        if ( {row,col} >= 038400 && {row,col} <= 038514) color_data <= 12'b111111110000; else
        if ( {row,col} >= 038515 && {row,col} <= 038895) color_data <= 12'b000010101110; else
        if ( {row,col} >= 038896 && {row,col} <= 038972) color_data <= 12'b111111111111; else
        if ( {row,col} >= 038973 && {row,col} <= 039039) color_data <= 12'b000010101110; else
        if ( {row,col} >= 039040 && {row,col} <= 039153) color_data <= 12'b111111110000; else
        if ( {row,col} >= 039154 && {row,col} <= 039536) color_data <= 12'b000010101110; else
        if ( {row,col} >= 039537 && {row,col} <= 039598) color_data <= 12'b111111111111; else
        if ( {row,col} >= 039599 && {row,col} <= 039602) color_data <= 12'b000010101110; else
        if ( {row,col} >= 039603 && {row,col} <= 039607) color_data <= 12'b111111111111; else
        if ( {row,col} >= 039608 && {row,col} <= 039679) color_data <= 12'b000010101110; else
        if ( {row,col} >= 039680 && {row,col} <= 039793) color_data <= 12'b111111110000; else
        if ( {row,col} >= 039794 && {row,col} <= 040182) color_data <= 12'b000010101110; else
        if ( {row,col} >= 040183 && {row,col} <= 040237) color_data <= 12'b111111111111; else
        if ( {row,col} >= 040238 && {row,col} <= 040319) color_data <= 12'b000010101110; else
        if ( {row,col} >= 040320 && {row,col} <= 040432) color_data <= 12'b111111110000; else
        if ( {row,col} >= 040433 && {row,col} <= 040827) color_data <= 12'b000010101110; else
        if ( {row,col} >= 040828 && {row,col} <= 040843) color_data <= 12'b111111111111; else
        if ( {row,col} >= 040844 && {row,col} <= 040844) color_data <= 12'b000010101110; else
        if ( {row,col} >= 040845 && {row,col} <= 040876) color_data <= 12'b111111111111; else
        if ( {row,col} >= 040877 && {row,col} <= 040959) color_data <= 12'b000010101110; else
        if ( {row,col} >= 040960 && {row,col} <= 041071) color_data <= 12'b111111110000; else
        if ( {row,col} >= 041072 && {row,col} <= 041469) color_data <= 12'b000010101110; else
        if ( {row,col} >= 041470 && {row,col} <= 041479) color_data <= 12'b111111111111; else
        if ( {row,col} >= 041480 && {row,col} <= 041485) color_data <= 12'b000010101110; else
        if ( {row,col} >= 041486 && {row,col} <= 041514) color_data <= 12'b111111111111; else
        if ( {row,col} >= 041515 && {row,col} <= 041599) color_data <= 12'b000010101110; else
        if ( {row,col} >= 041600 && {row,col} <= 041711) color_data <= 12'b111111110000; else
        if ( {row,col} >= 041712 && {row,col} <= 042127) color_data <= 12'b000010101110; else
        if ( {row,col} >= 042128 && {row,col} <= 042152) color_data <= 12'b111111111111; else
        if ( {row,col} >= 042153 && {row,col} <= 042239) color_data <= 12'b000010101110; else
        if ( {row,col} >= 042240 && {row,col} <= 042350) color_data <= 12'b111111110000; else
        if ( {row,col} >= 042351 && {row,col} <= 042770) color_data <= 12'b000010101110; else
        if ( {row,col} >= 042771 && {row,col} <= 042790) color_data <= 12'b111111111111; else
        if ( {row,col} >= 042791 && {row,col} <= 042879) color_data <= 12'b000010101110; else
        if ( {row,col} >= 042880 && {row,col} <= 042989) color_data <= 12'b111111110000; else
        if ( {row,col} >= 042990 && {row,col} <= 043414) color_data <= 12'b000010101110; else
        if ( {row,col} >= 043415 && {row,col} <= 043426) color_data <= 12'b111111111111; else
        if ( {row,col} >= 043427 && {row,col} <= 043519) color_data <= 12'b000010101110; else
        if ( {row,col} >= 043520 && {row,col} <= 043629) color_data <= 12'b111111110000; else
        if ( {row,col} >= 043630 && {row,col} <= 044159) color_data <= 12'b000010101110; else
        if ( {row,col} >= 044160 && {row,col} <= 044268) color_data <= 12'b111111110000; else
        if ( {row,col} >= 044269 && {row,col} <= 044799) color_data <= 12'b000010101110; else
        if ( {row,col} >= 044800 && {row,col} <= 044907) color_data <= 12'b111111110000; else
        if ( {row,col} >= 044908 && {row,col} <= 045439) color_data <= 12'b000010101110; else
        if ( {row,col} >= 045440 && {row,col} <= 045546) color_data <= 12'b111111110000; else
        if ( {row,col} >= 045547 && {row,col} <= 046079) color_data <= 12'b000010101110; else
        if ( {row,col} >= 046080 && {row,col} <= 046185) color_data <= 12'b111111110000; else
        if ( {row,col} >= 046186 && {row,col} <= 046719) color_data <= 12'b000010101110; else
        if ( {row,col} >= 046720 && {row,col} <= 046825) color_data <= 12'b111111110000; else
        if ( {row,col} >= 046826 && {row,col} <= 047359) color_data <= 12'b000010101110; else
        if ( {row,col} >= 047360 && {row,col} <= 047464) color_data <= 12'b111111110000; else
        if ( {row,col} >= 047465 && {row,col} <= 047999) color_data <= 12'b000010101110; else
        if ( {row,col} >= 048000 && {row,col} <= 048103) color_data <= 12'b111111110000; else
        if ( {row,col} >= 048104 && {row,col} <= 048639) color_data <= 12'b000010101110; else
        if ( {row,col} >= 048640 && {row,col} <= 048742) color_data <= 12'b111111110000; else
        if ( {row,col} >= 048743 && {row,col} <= 049279) color_data <= 12'b000010101110; else
        if ( {row,col} >= 049280 && {row,col} <= 049381) color_data <= 12'b111111110000; else
        if ( {row,col} >= 049382 && {row,col} <= 049919) color_data <= 12'b000010101110; else
        if ( {row,col} >= 049920 && {row,col} <= 050020) color_data <= 12'b111111110000; else
        if ( {row,col} >= 050021 && {row,col} <= 050559) color_data <= 12'b000010101110; else
        if ( {row,col} >= 050560 && {row,col} <= 050659) color_data <= 12'b111111110000; else
        if ( {row,col} >= 050660 && {row,col} <= 051199) color_data <= 12'b000010101110; else
        if ( {row,col} >= 051200 && {row,col} <= 051298) color_data <= 12'b111111110000; else
        if ( {row,col} >= 051299 && {row,col} <= 051839) color_data <= 12'b000010101110; else
        if ( {row,col} >= 051840 && {row,col} <= 051937) color_data <= 12'b111111110000; else
        if ( {row,col} >= 051938 && {row,col} <= 052479) color_data <= 12'b000010101110; else
        if ( {row,col} >= 052480 && {row,col} <= 052576) color_data <= 12'b111111110000; else
        if ( {row,col} >= 052577 && {row,col} <= 053119) color_data <= 12'b000010101110; else
        if ( {row,col} >= 053120 && {row,col} <= 053215) color_data <= 12'b111111110000; else
        if ( {row,col} >= 053216 && {row,col} <= 053759) color_data <= 12'b000010101110; else
        if ( {row,col} >= 053760 && {row,col} <= 053854) color_data <= 12'b111111110000; else
        if ( {row,col} >= 053855 && {row,col} <= 054399) color_data <= 12'b000010101110; else
        if ( {row,col} >= 054400 && {row,col} <= 054493) color_data <= 12'b111111110000; else
        if ( {row,col} >= 054494 && {row,col} <= 055039) color_data <= 12'b000010101110; else
        if ( {row,col} >= 055040 && {row,col} <= 055132) color_data <= 12'b111111110000; else
        if ( {row,col} >= 055133 && {row,col} <= 055679) color_data <= 12'b000010101110; else
        if ( {row,col} >= 055680 && {row,col} <= 055771) color_data <= 12'b111111110000; else
        if ( {row,col} >= 055772 && {row,col} <= 056319) color_data <= 12'b000010101110; else
        if ( {row,col} >= 056320 && {row,col} <= 056410) color_data <= 12'b111111110000; else
        if ( {row,col} >= 056411 && {row,col} <= 056959) color_data <= 12'b000010101110; else
        if ( {row,col} >= 056960 && {row,col} <= 057049) color_data <= 12'b111111110000; else
        if ( {row,col} >= 057050 && {row,col} <= 057599) color_data <= 12'b000010101110; else
        if ( {row,col} >= 057600 && {row,col} <= 057688) color_data <= 12'b111111110000; else
        if ( {row,col} >= 057689 && {row,col} <= 058239) color_data <= 12'b000010101110; else
        if ( {row,col} >= 058240 && {row,col} <= 058326) color_data <= 12'b111111110000; else
        if ( {row,col} >= 058327 && {row,col} <= 058879) color_data <= 12'b000010101110; else
        if ( {row,col} >= 058880 && {row,col} <= 058965) color_data <= 12'b111111110000; else
        if ( {row,col} >= 058966 && {row,col} <= 059519) color_data <= 12'b000010101110; else
        if ( {row,col} >= 059520 && {row,col} <= 059604) color_data <= 12'b111111110000; else
        if ( {row,col} >= 059605 && {row,col} <= 060159) color_data <= 12'b000010101110; else
        if ( {row,col} >= 060160 && {row,col} <= 060243) color_data <= 12'b111111110000; else
        if ( {row,col} >= 060244 && {row,col} <= 060799) color_data <= 12'b000010101110; else
        if ( {row,col} >= 060800 && {row,col} <= 060881) color_data <= 12'b111111110000; else
        if ( {row,col} >= 060882 && {row,col} <= 061439) color_data <= 12'b000010101110; else
        if ( {row,col} >= 061440 && {row,col} <= 061520) color_data <= 12'b111111110000; else
        if ( {row,col} >= 061521 && {row,col} <= 062079) color_data <= 12'b000010101110; else
        if ( {row,col} >= 062080 && {row,col} <= 062158) color_data <= 12'b111111110000; else
        if ( {row,col} >= 062159 && {row,col} <= 062719) color_data <= 12'b000010101110; else
        if ( {row,col} >= 062720 && {row,col} <= 062797) color_data <= 12'b111111110000; else
        if ( {row,col} >= 062798 && {row,col} <= 063359) color_data <= 12'b000010101110; else
        if ( {row,col} >= 063360 && {row,col} <= 063436) color_data <= 12'b111111110000; else
        if ( {row,col} >= 063437 && {row,col} <= 063999) color_data <= 12'b000010101110; else
        if ( {row,col} >= 064000 && {row,col} <= 064074) color_data <= 12'b111111110000; else
        if ( {row,col} >= 064075 && {row,col} <= 064639) color_data <= 12'b000010101110; else
        if ( {row,col} >= 064640 && {row,col} <= 064713) color_data <= 12'b111111110000; else
        if ( {row,col} >= 064714 && {row,col} <= 065279) color_data <= 12'b000010101110; else
        if ( {row,col} >= 065280 && {row,col} <= 065351) color_data <= 12'b111111110000; else
        if ( {row,col} >= 065352 && {row,col} <= 065919) color_data <= 12'b000010101110; else
        if ( {row,col} >= 065920 && {row,col} <= 065989) color_data <= 12'b111111110000; else
        if ( {row,col} >= 065990 && {row,col} <= 066559) color_data <= 12'b000010101110; else
        if ( {row,col} >= 066560 && {row,col} <= 066627) color_data <= 12'b111111110000; else
        if ( {row,col} >= 066628 && {row,col} <= 067199) color_data <= 12'b000010101110; else
        if ( {row,col} >= 067200 && {row,col} <= 067265) color_data <= 12'b111111110000; else
        if ( {row,col} >= 067266 && {row,col} <= 067839) color_data <= 12'b000010101110; else
        if ( {row,col} >= 067840 && {row,col} <= 067904) color_data <= 12'b111111110000; else
        if ( {row,col} >= 067905 && {row,col} <= 068479) color_data <= 12'b000010101110; else
        if ( {row,col} >= 068480 && {row,col} <= 068542) color_data <= 12'b111111110000; else
        if ( {row,col} >= 068543 && {row,col} <= 069119) color_data <= 12'b000010101110; else
        if ( {row,col} >= 069120 && {row,col} <= 069180) color_data <= 12'b111111110000; else
        if ( {row,col} >= 069181 && {row,col} <= 069759) color_data <= 12'b000010101110; else
        if ( {row,col} >= 069760 && {row,col} <= 069817) color_data <= 12'b111111110000; else
        if ( {row,col} >= 069818 && {row,col} <= 070399) color_data <= 12'b000010101110; else
        if ( {row,col} >= 070400 && {row,col} <= 070455) color_data <= 12'b111111110000; else
        if ( {row,col} >= 070456 && {row,col} <= 071039) color_data <= 12'b000010101110; else
        if ( {row,col} >= 071040 && {row,col} <= 071093) color_data <= 12'b111111110000; else
        if ( {row,col} >= 071094 && {row,col} <= 071679) color_data <= 12'b000010101110; else
        if ( {row,col} >= 071680 && {row,col} <= 071731) color_data <= 12'b111111110000; else
        if ( {row,col} >= 071732 && {row,col} <= 072319) color_data <= 12'b000010101110; else
        if ( {row,col} >= 072320 && {row,col} <= 072368) color_data <= 12'b111111110000; else
        if ( {row,col} >= 072369 && {row,col} <= 072959) color_data <= 12'b000010101110; else
        if ( {row,col} >= 072960 && {row,col} <= 073005) color_data <= 12'b111111110000; else
        if ( {row,col} >= 073006 && {row,col} <= 073599) color_data <= 12'b000010101110; else
        if ( {row,col} >= 073600 && {row,col} <= 073642) color_data <= 12'b111111110000; else
        if ( {row,col} >= 073643 && {row,col} <= 074239) color_data <= 12'b000010101110; else
        if ( {row,col} >= 074240 && {row,col} <= 074279) color_data <= 12'b111111110000; else
        if ( {row,col} >= 074280 && {row,col} <= 074879) color_data <= 12'b000010101110; else
        if ( {row,col} >= 074880 && {row,col} <= 074914) color_data <= 12'b111111110000; else
        if ( {row,col} >= 074915 && {row,col} <= 075519) color_data <= 12'b000010101110; else
        if ( {row,col} >= 075520 && {row,col} <= 075550) color_data <= 12'b111111110000; else
        if ( {row,col} >= 075551 && {row,col} <= 076159) color_data <= 12'b000010101110; else
        if ( {row,col} >= 076160 && {row,col} <= 076186) color_data <= 12'b111111110000; else
        if ( {row,col} >= 076187 && {row,col} <= 076799) color_data <= 12'b000010101110; else
        if ( {row,col} >= 076800 && {row,col} <= 076819) color_data <= 12'b111111110000; else
        if ( {row,col} >= 076820 && {row,col} <= 077439) color_data <= 12'b000010101110; else
        if ( {row,col} >= 077440 && {row,col} <= 077450) color_data <= 12'b111111110000; else
        if ( {row,col} >= 077451 && {row,col} <= 202879) color_data <= 12'b000010101110; else
        if ( {row,col} >= 202880 && {row,col} <= 226559) color_data <= 12'b001010110100; else
        if ( {row,col} >= 226560 && {row,col} <= 249364) color_data <= 12'b000000000000; else
        if ( {row,col} >= 249365 && {row,col} <= 249407) color_data <= 12'b111111110000; else
        if ( {row,col} >= 249408 && {row,col} <= 249515) color_data <= 12'b000000000000; else
        if ( {row,col} >= 249516 && {row,col} <= 249558) color_data <= 12'b111111110000; else
        if ( {row,col} >= 249559 && {row,col} <= 249927) color_data <= 12'b000000000000; else
        if ( {row,col} >= 249928 && {row,col} <= 249970) color_data <= 12'b111111110000; else
        if ( {row,col} >= 249971 && {row,col} <= 250004) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250005 && {row,col} <= 250047) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250048 && {row,col} <= 250083) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250084 && {row,col} <= 250126) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250127 && {row,col} <= 250155) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250156 && {row,col} <= 250198) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250199 && {row,col} <= 250266) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250267 && {row,col} <= 250309) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250310 && {row,col} <= 250337) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250338 && {row,col} <= 250380) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250381 && {row,col} <= 250485) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250486 && {row,col} <= 250528) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250529 && {row,col} <= 250567) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250568 && {row,col} <= 250610) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250611 && {row,col} <= 250644) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250645 && {row,col} <= 250687) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250688 && {row,col} <= 250723) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250724 && {row,col} <= 250766) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250767 && {row,col} <= 250795) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250796 && {row,col} <= 250838) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250839 && {row,col} <= 250906) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250907 && {row,col} <= 250949) color_data <= 12'b111111110000; else
        if ( {row,col} >= 250950 && {row,col} <= 250977) color_data <= 12'b000000000000; else
        if ( {row,col} >= 250978 && {row,col} <= 251020) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251021 && {row,col} <= 251050) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251051 && {row,col} <= 251093) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251094 && {row,col} <= 251125) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251126 && {row,col} <= 251168) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251169 && {row,col} <= 251207) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251208 && {row,col} <= 251250) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251251 && {row,col} <= 251284) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251285 && {row,col} <= 251327) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251328 && {row,col} <= 251363) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251364 && {row,col} <= 251406) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251407 && {row,col} <= 251435) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251436 && {row,col} <= 251478) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251479 && {row,col} <= 251546) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251547 && {row,col} <= 251589) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251590 && {row,col} <= 251617) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251618 && {row,col} <= 251660) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251661 && {row,col} <= 251690) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251691 && {row,col} <= 251733) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251734 && {row,col} <= 251765) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251766 && {row,col} <= 251808) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251809 && {row,col} <= 251847) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251848 && {row,col} <= 251890) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251891 && {row,col} <= 251924) color_data <= 12'b000000000000; else
        if ( {row,col} >= 251925 && {row,col} <= 251967) color_data <= 12'b111111110000; else
        if ( {row,col} >= 251968 && {row,col} <= 252003) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252004 && {row,col} <= 252046) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252047 && {row,col} <= 252075) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252076 && {row,col} <= 252118) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252119 && {row,col} <= 252186) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252187 && {row,col} <= 252229) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252230 && {row,col} <= 252257) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252258 && {row,col} <= 252300) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252301 && {row,col} <= 252330) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252331 && {row,col} <= 252373) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252374 && {row,col} <= 252405) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252406 && {row,col} <= 252448) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252449 && {row,col} <= 252487) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252488 && {row,col} <= 252530) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252531 && {row,col} <= 252564) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252565 && {row,col} <= 252607) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252608 && {row,col} <= 252643) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252644 && {row,col} <= 252686) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252687 && {row,col} <= 252715) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252716 && {row,col} <= 252758) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252759 && {row,col} <= 252826) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252827 && {row,col} <= 252869) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252870 && {row,col} <= 252897) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252898 && {row,col} <= 252940) color_data <= 12'b111111110000; else
        if ( {row,col} >= 252941 && {row,col} <= 252970) color_data <= 12'b000000000000; else
        if ( {row,col} >= 252971 && {row,col} <= 253013) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253014 && {row,col} <= 253045) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253046 && {row,col} <= 253088) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253089 && {row,col} <= 253127) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253128 && {row,col} <= 253170) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253171 && {row,col} <= 253204) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253205 && {row,col} <= 253247) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253248 && {row,col} <= 253283) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253284 && {row,col} <= 253326) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253327 && {row,col} <= 253355) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253356 && {row,col} <= 253398) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253399 && {row,col} <= 253466) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253467 && {row,col} <= 253509) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253510 && {row,col} <= 253537) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253538 && {row,col} <= 253580) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253581 && {row,col} <= 253610) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253611 && {row,col} <= 253653) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253654 && {row,col} <= 253685) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253686 && {row,col} <= 253728) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253729 && {row,col} <= 253767) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253768 && {row,col} <= 253810) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253811 && {row,col} <= 253844) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253845 && {row,col} <= 253887) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253888 && {row,col} <= 253923) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253924 && {row,col} <= 253966) color_data <= 12'b111111110000; else
        if ( {row,col} >= 253967 && {row,col} <= 253995) color_data <= 12'b000000000000; else
        if ( {row,col} >= 253996 && {row,col} <= 254038) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254039 && {row,col} <= 254106) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254107 && {row,col} <= 254149) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254150 && {row,col} <= 254177) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254178 && {row,col} <= 254220) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254221 && {row,col} <= 254250) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254251 && {row,col} <= 254293) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254294 && {row,col} <= 254325) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254326 && {row,col} <= 254368) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254369 && {row,col} <= 254407) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254408 && {row,col} <= 254450) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254451 && {row,col} <= 254484) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254485 && {row,col} <= 254527) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254528 && {row,col} <= 254563) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254564 && {row,col} <= 254606) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254607 && {row,col} <= 254635) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254636 && {row,col} <= 254678) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254679 && {row,col} <= 254746) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254747 && {row,col} <= 254789) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254790 && {row,col} <= 254817) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254818 && {row,col} <= 254860) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254861 && {row,col} <= 254890) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254891 && {row,col} <= 254933) color_data <= 12'b111111110000; else
        if ( {row,col} >= 254934 && {row,col} <= 254965) color_data <= 12'b000000000000; else
        if ( {row,col} >= 254966 && {row,col} <= 255008) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255009 && {row,col} <= 255047) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255048 && {row,col} <= 255090) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255091 && {row,col} <= 255124) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255125 && {row,col} <= 255167) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255168 && {row,col} <= 255203) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255204 && {row,col} <= 255246) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255247 && {row,col} <= 255275) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255276 && {row,col} <= 255318) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255319 && {row,col} <= 255386) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255387 && {row,col} <= 255429) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255430 && {row,col} <= 255457) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255458 && {row,col} <= 255500) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255501 && {row,col} <= 255530) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255531 && {row,col} <= 255573) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255574 && {row,col} <= 255605) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255606 && {row,col} <= 255648) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255649 && {row,col} <= 255687) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255688 && {row,col} <= 255730) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255731 && {row,col} <= 255764) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255765 && {row,col} <= 255807) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255808 && {row,col} <= 255843) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255844 && {row,col} <= 255886) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255887 && {row,col} <= 255915) color_data <= 12'b000000000000; else
        if ( {row,col} >= 255916 && {row,col} <= 255958) color_data <= 12'b111111110000; else
        if ( {row,col} >= 255959 && {row,col} <= 256026) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256027 && {row,col} <= 256069) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256070 && {row,col} <= 256097) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256098 && {row,col} <= 256140) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256141 && {row,col} <= 256170) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256171 && {row,col} <= 256213) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256214 && {row,col} <= 256245) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256246 && {row,col} <= 256288) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256289 && {row,col} <= 256327) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256328 && {row,col} <= 256370) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256371 && {row,col} <= 256483) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256484 && {row,col} <= 256526) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256527 && {row,col} <= 256666) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256667 && {row,col} <= 256709) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256710 && {row,col} <= 256737) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256738 && {row,col} <= 256780) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256781 && {row,col} <= 256810) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256811 && {row,col} <= 256853) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256854 && {row,col} <= 256885) color_data <= 12'b000000000000; else
        if ( {row,col} >= 256886 && {row,col} <= 256928) color_data <= 12'b111111110000; else
        if ( {row,col} >= 256929 && {row,col} <= 257450) color_data <= 12'b000000000000; else
        if ( {row,col} >= 257451 && {row,col} <= 257493) color_data <= 12'b111111110000; else
        if ( {row,col} >= 257494 && {row,col} <= 279679) color_data <= 12'b000000000000; else
        if ( {row,col} >= 279680 && {row,col} < 307200) color_data <= 12'b001010110100; else
        // default case
        color_data <= 12'b000000000000;
    end
endmodule
