module nine_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "distributed" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		10'b0000101010: color_data = 12'b000000000000;
		10'b0000101011: color_data = 12'b000000000000;
		10'b0000101100: color_data = 12'b000000000000;
		10'b0000101101: color_data = 12'b000000000000;
		10'b0000101110: color_data = 12'b000000000000;
		10'b0001001000: color_data = 12'b000000000000;
		10'b0001001001: color_data = 12'b000000000000;
		10'b0001001010: color_data = 12'b000000000000;
		10'b0001001011: color_data = 12'b000000000000;
		10'b0001001100: color_data = 12'b000000000000;
		10'b0001001101: color_data = 12'b000000000000;
		10'b0001001110: color_data = 12'b000000000000;
		10'b0001001111: color_data = 12'b000000000000;
		10'b0001100110: color_data = 12'b000000000000;
		10'b0001100111: color_data = 12'b000000000000;
		10'b0001101000: color_data = 12'b000000000000;
		10'b0001101001: color_data = 12'b000000000000;
		10'b0001101010: color_data = 12'b000000000000;
		10'b0001101011: color_data = 12'b000000000000;
		10'b0001101100: color_data = 12'b000000000000;
		10'b0001101101: color_data = 12'b000000000000;
		10'b0001101110: color_data = 12'b000000000000;
		10'b0001101111: color_data = 12'b000000000000;
		10'b0001110000: color_data = 12'b000000000000;
		10'b0001110001: color_data = 12'b000000000000;
		10'b0010000110: color_data = 12'b000000000000;
		10'b0010000111: color_data = 12'b000000000000;
		10'b0010001000: color_data = 12'b000000000000;
		10'b0010001001: color_data = 12'b000000000000;
		10'b0010001110: color_data = 12'b000000000000;
		10'b0010001111: color_data = 12'b000000000000;
		10'b0010010000: color_data = 12'b000000000000;
		10'b0010010001: color_data = 12'b000000000000;
		10'b0010010010: color_data = 12'b000000000000;
		10'b0010010011: color_data = 12'b000000000000;
		10'b0010100101: color_data = 12'b000000000000;
		10'b0010100110: color_data = 12'b000000000000;
		10'b0010100111: color_data = 12'b000000000000;
		10'b0010101000: color_data = 12'b000000000000;
		10'b0010101111: color_data = 12'b000000000000;
		10'b0010110000: color_data = 12'b000000000000;
		10'b0010110001: color_data = 12'b000000000000;
		10'b0010110010: color_data = 12'b000000000000;
		10'b0010110011: color_data = 12'b000000000000;
		10'b0011000101: color_data = 12'b000000000000;
		10'b0011000110: color_data = 12'b000000000000;
		10'b0011000111: color_data = 12'b000000000000;
		10'b0011010000: color_data = 12'b000000000000;
		10'b0011010001: color_data = 12'b000000000000;
		10'b0011010010: color_data = 12'b000000000000;
		10'b0011010011: color_data = 12'b000000000000;
		10'b0011100100: color_data = 12'b000000000000;
		10'b0011100101: color_data = 12'b000000000000;
		10'b0011100110: color_data = 12'b000000000000;
		10'b0011110001: color_data = 12'b000000000000;
		10'b0011110010: color_data = 12'b000000000000;
		10'b0011110011: color_data = 12'b000000000000;
		10'b0100000100: color_data = 12'b000000000000;
		10'b0100000101: color_data = 12'b000000000000;
		10'b0100000110: color_data = 12'b000000000000;
		10'b0100010001: color_data = 12'b000000000000;
		10'b0100010010: color_data = 12'b000000000000;
		10'b0100010011: color_data = 12'b000000000000;
		10'b0100100100: color_data = 12'b000000000000;
		10'b0100100101: color_data = 12'b000000000000;
		10'b0100100110: color_data = 12'b000000000000;
		10'b0100110001: color_data = 12'b000000000000;
		10'b0100110010: color_data = 12'b000000000000;
		10'b0100110011: color_data = 12'b000000000000;
		10'b0101000100: color_data = 12'b000000000000;
		10'b0101000101: color_data = 12'b000000000000;
		10'b0101000110: color_data = 12'b000000000000;
		10'b0101010001: color_data = 12'b000000000000;
		10'b0101010010: color_data = 12'b000000000000;
		10'b0101010011: color_data = 12'b000000000000;
		10'b0101100100: color_data = 12'b000000000000;
		10'b0101100101: color_data = 12'b000000000000;
		10'b0101100110: color_data = 12'b000000000000;
		10'b0101100111: color_data = 12'b000000000000;
		10'b0101110000: color_data = 12'b000000000000;
		10'b0101110001: color_data = 12'b000000000000;
		10'b0101110010: color_data = 12'b000000000000;
		10'b0101110011: color_data = 12'b000000000000;
		10'b0110000101: color_data = 12'b000000000000;
		10'b0110000110: color_data = 12'b000000000000;
		10'b0110000111: color_data = 12'b000000000000;
		10'b0110010000: color_data = 12'b000000000000;
		10'b0110010001: color_data = 12'b000000000000;
		10'b0110010010: color_data = 12'b000000000000;
		10'b0110010011: color_data = 12'b000000000000;
		10'b0110100110: color_data = 12'b000000000000;
		10'b0110100111: color_data = 12'b000000000000;
		10'b0110101000: color_data = 12'b000000000000;
		10'b0110101001: color_data = 12'b000000000000;
		10'b0110101110: color_data = 12'b000000000000;
		10'b0110101111: color_data = 12'b000000000000;
		10'b0110110000: color_data = 12'b000000000000;
		10'b0110110001: color_data = 12'b000000000000;
		10'b0110110010: color_data = 12'b000000000000;
		10'b0110110011: color_data = 12'b000000000000;
		10'b0111000110: color_data = 12'b000000000000;
		10'b0111000111: color_data = 12'b000000000000;
		10'b0111001000: color_data = 12'b000000000000;
		10'b0111001001: color_data = 12'b000000000000;
		10'b0111001010: color_data = 12'b000000000000;
		10'b0111001011: color_data = 12'b000000000000;
		10'b0111001100: color_data = 12'b000000000000;
		10'b0111001101: color_data = 12'b000000000000;
		10'b0111001110: color_data = 12'b000000000000;
		10'b0111001111: color_data = 12'b000000000000;
		10'b0111010000: color_data = 12'b000000000000;
		10'b0111010001: color_data = 12'b000000000000;
		10'b0111010010: color_data = 12'b000000000000;
		10'b0111010011: color_data = 12'b000000000000;
		10'b0111101000: color_data = 12'b000000000000;
		10'b0111101001: color_data = 12'b000000000000;
		10'b0111101010: color_data = 12'b000000000000;
		10'b0111101011: color_data = 12'b000000000000;
		10'b0111101100: color_data = 12'b000000000000;
		10'b0111101101: color_data = 12'b000000000000;
		10'b0111101110: color_data = 12'b000000000000;
		10'b0111101111: color_data = 12'b000000000000;
		10'b0111110000: color_data = 12'b000000000000;
		10'b0111110001: color_data = 12'b000000000000;
		10'b0111110010: color_data = 12'b000000000000;
		10'b0111110011: color_data = 12'b000000000000;
		10'b1000001001: color_data = 12'b000000000000;
		10'b1000001010: color_data = 12'b000000000000;
		10'b1000001011: color_data = 12'b000000000000;
		10'b1000001100: color_data = 12'b000000000000;
		10'b1000001101: color_data = 12'b000000000000;
		10'b1000001110: color_data = 12'b000000000000;
		10'b1000010001: color_data = 12'b000000000000;
		10'b1000010010: color_data = 12'b000000000000;
		10'b1000010011: color_data = 12'b000000000000;
		10'b1000110001: color_data = 12'b000000000000;
		10'b1000110010: color_data = 12'b000000000000;
		10'b1000110011: color_data = 12'b000000000000;
		10'b1001010001: color_data = 12'b000000000000;
		10'b1001010010: color_data = 12'b000000000000;
		10'b1001010011: color_data = 12'b000000000000;
		10'b1001110001: color_data = 12'b000000000000;
		10'b1001110010: color_data = 12'b000000000000;
		10'b1001110011: color_data = 12'b000000000000;
		10'b1010010001: color_data = 12'b000000000000;
		10'b1010010010: color_data = 12'b000000000000;
		10'b1010010011: color_data = 12'b000000000000;
		10'b1010110001: color_data = 12'b000000000000;
		10'b1010110010: color_data = 12'b000000000000;
		10'b1010110011: color_data = 12'b000000000000;
		10'b1011010001: color_data = 12'b000000000000;
		10'b1011010010: color_data = 12'b000000000000;
		10'b1011010011: color_data = 12'b000000000000;
		10'b1011110001: color_data = 12'b000000000000;
		10'b1011110010: color_data = 12'b000000000000;
		10'b1011110011: color_data = 12'b000000000000;
		10'b1100010001: color_data = 12'b000000000000;
		10'b1100010010: color_data = 12'b000000000000;
		10'b1100010011: color_data = 12'b000000000000;
		10'b1100110001: color_data = 12'b000000000000;
		10'b1100110010: color_data = 12'b000000000000;
		10'b1100110011: color_data = 12'b000000000000;
		10'b1101010001: color_data = 12'b000000000000;
		10'b1101010010: color_data = 12'b000000000000;
		10'b1101010011: color_data = 12'b000000000000;
		10'b1101110001: color_data = 12'b000000000000;
		10'b1101110010: color_data = 12'b000000000000;
		10'b1101110011: color_data = 12'b000000000000;
		10'b1110010001: color_data = 12'b000000000000;
		10'b1110010010: color_data = 12'b000000000000;
		10'b1110010011: color_data = 12'b000000000000;
        default: color_data = 12'b111111111111;
	endcase
endmodule