`timescale 1ns / 1ps
module background_rom (
    input wire clk,
    input wire [8:0] row,
    input wire [9:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 640 + col) >= 0 && (row * 640 + col) <= 131) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 132 && (row * 640 + col) <= 639) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 640 && (row * 640 + col) <= 771) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 772 && (row * 640 + col) <= 1279) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 1280 && (row * 640 + col) <= 1411) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 1412 && (row * 640 + col) <= 1919) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 1920 && (row * 640 + col) <= 2051) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 2052 && (row * 640 + col) <= 2559) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 2560 && (row * 640 + col) <= 2691) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 2692 && (row * 640 + col) <= 3199) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 3200 && (row * 640 + col) <= 3331) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 3332 && (row * 640 + col) <= 3839) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 3840 && (row * 640 + col) <= 3971) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 3972 && (row * 640 + col) <= 4479) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 4480 && (row * 640 + col) <= 4611) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 4612 && (row * 640 + col) <= 5119) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 5120 && (row * 640 + col) <= 5251) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 5252 && (row * 640 + col) <= 5759) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 5760 && (row * 640 + col) <= 5890) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 5891 && (row * 640 + col) <= 6399) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 6400 && (row * 640 + col) <= 6530) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 6531 && (row * 640 + col) <= 7039) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 7040 && (row * 640 + col) <= 7170) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 7171 && (row * 640 + col) <= 7679) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 7680 && (row * 640 + col) <= 7810) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 7811 && (row * 640 + col) <= 8319) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 8320 && (row * 640 + col) <= 8450) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 8451 && (row * 640 + col) <= 8959) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 8960 && (row * 640 + col) <= 9090) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 9091 && (row * 640 + col) <= 9507) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 9508 && (row * 640 + col) <= 9514) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 9515 && (row * 640 + col) <= 9525) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 9526 && (row * 640 + col) <= 9533) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 9534 && (row * 640 + col) <= 9599) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 9600 && (row * 640 + col) <= 9730) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 9731 && (row * 640 + col) <= 10143) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 10144 && (row * 640 + col) <= 10157) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 10158 && (row * 640 + col) <= 10162) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 10163 && (row * 640 + col) <= 10177) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 10178 && (row * 640 + col) <= 10239) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 10240 && (row * 640 + col) <= 10370) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 10371 && (row * 640 + col) <= 10765) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 10766 && (row * 640 + col) <= 10776) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 10777 && (row * 640 + col) <= 10781) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 10782 && (row * 640 + col) <= 10819) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 10820 && (row * 640 + col) <= 10879) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 10880 && (row * 640 + col) <= 11010) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 11011 && (row * 640 + col) <= 11402) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 11403 && (row * 640 + col) <= 11461) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 11462 && (row * 640 + col) <= 11519) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 11520 && (row * 640 + col) <= 11649) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 11650 && (row * 640 + col) <= 12040) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 12041 && (row * 640 + col) <= 12102) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 12103 && (row * 640 + col) <= 12159) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 12160 && (row * 640 + col) <= 12289) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 12290 && (row * 640 + col) <= 12662) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 12663 && (row * 640 + col) <= 12676) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 12677 && (row * 640 + col) <= 12678) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 12679 && (row * 640 + col) <= 12743) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 12744 && (row * 640 + col) <= 12799) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 12800 && (row * 640 + col) <= 12929) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 12930 && (row * 640 + col) <= 13299) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 13300 && (row * 640 + col) <= 13384) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 13385 && (row * 640 + col) <= 13439) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 13440 && (row * 640 + col) <= 13569) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 13570 && (row * 640 + col) <= 13937) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 13938 && (row * 640 + col) <= 14026) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 14027 && (row * 640 + col) <= 14079) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 14080 && (row * 640 + col) <= 14209) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 14210 && (row * 640 + col) <= 14575) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 14576 && (row * 640 + col) <= 14668) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 14669 && (row * 640 + col) <= 14719) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 14720 && (row * 640 + col) <= 14849) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 14850 && (row * 640 + col) <= 15214) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 15215 && (row * 640 + col) <= 15310) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 15311 && (row * 640 + col) <= 15359) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 15360 && (row * 640 + col) <= 15488) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 15489 && (row * 640 + col) <= 15853) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 15854 && (row * 640 + col) <= 15951) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 15952 && (row * 640 + col) <= 15999) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 16000 && (row * 640 + col) <= 16128) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 16129 && (row * 640 + col) <= 16492) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 16493 && (row * 640 + col) <= 16592) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 16593 && (row * 640 + col) <= 16639) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 16640 && (row * 640 + col) <= 16768) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 16769 && (row * 640 + col) <= 17131) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 17132 && (row * 640 + col) <= 17233) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17234 && (row * 640 + col) <= 17279) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 17280 && (row * 640 + col) <= 17408) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 17409 && (row * 640 + col) <= 17771) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 17772 && (row * 640 + col) <= 17874) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 17875 && (row * 640 + col) <= 17919) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 17920 && (row * 640 + col) <= 18047) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 18048 && (row * 640 + col) <= 18410) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 18411 && (row * 640 + col) <= 18514) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 18515 && (row * 640 + col) <= 18559) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 18560 && (row * 640 + col) <= 18687) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 18688 && (row * 640 + col) <= 19050) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 19051 && (row * 640 + col) <= 19154) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19155 && (row * 640 + col) <= 19199) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 19200 && (row * 640 + col) <= 19327) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 19328 && (row * 640 + col) <= 19690) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 19691 && (row * 640 + col) <= 19795) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 19796 && (row * 640 + col) <= 19839) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 19840 && (row * 640 + col) <= 19967) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 19968 && (row * 640 + col) <= 20326) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 20327 && (row * 640 + col) <= 20435) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 20436 && (row * 640 + col) <= 20479) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 20480 && (row * 640 + col) <= 20606) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 20607 && (row * 640 + col) <= 20964) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 20965 && (row * 640 + col) <= 21074) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21075 && (row * 640 + col) <= 21119) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 21120 && (row * 640 + col) <= 21246) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 21247 && (row * 640 + col) <= 21602) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 21603 && (row * 640 + col) <= 21714) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 21715 && (row * 640 + col) <= 21759) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 21760 && (row * 640 + col) <= 21886) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 21887 && (row * 640 + col) <= 22240) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 22241 && (row * 640 + col) <= 22355) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22356 && (row * 640 + col) <= 22399) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 22400 && (row * 640 + col) <= 22525) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 22526 && (row * 640 + col) <= 22880) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 22881 && (row * 640 + col) <= 22995) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 22996 && (row * 640 + col) <= 23039) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 23040 && (row * 640 + col) <= 23165) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 23166 && (row * 640 + col) <= 23519) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 23520 && (row * 640 + col) <= 23636) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 23637 && (row * 640 + col) <= 23679) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 23680 && (row * 640 + col) <= 23805) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 23806 && (row * 640 + col) <= 24158) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 24159 && (row * 640 + col) <= 24276) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24277 && (row * 640 + col) <= 24319) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 24320 && (row * 640 + col) <= 24444) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 24445 && (row * 640 + col) <= 24798) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 24799 && (row * 640 + col) <= 24917) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 24918 && (row * 640 + col) <= 24959) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 24960 && (row * 640 + col) <= 25084) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 25085 && (row * 640 + col) <= 25438) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 25439 && (row * 640 + col) <= 25557) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 25558 && (row * 640 + col) <= 25599) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 25600 && (row * 640 + col) <= 25724) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 25725 && (row * 640 + col) <= 26078) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 26079 && (row * 640 + col) <= 26197) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26198 && (row * 640 + col) <= 26239) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 26240 && (row * 640 + col) <= 26363) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 26364 && (row * 640 + col) <= 26718) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 26719 && (row * 640 + col) <= 26837) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 26838 && (row * 640 + col) <= 26879) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 26880 && (row * 640 + col) <= 27003) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 27004 && (row * 640 + col) <= 27359) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 27360 && (row * 640 + col) <= 27477) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 27478 && (row * 640 + col) <= 27519) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 27520 && (row * 640 + col) <= 27642) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 27643 && (row * 640 + col) <= 27999) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 28000 && (row * 640 + col) <= 28116) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28117 && (row * 640 + col) <= 28159) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 28160 && (row * 640 + col) <= 28282) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 28283 && (row * 640 + col) <= 28640) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 28641 && (row * 640 + col) <= 28756) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 28757 && (row * 640 + col) <= 28799) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 28800 && (row * 640 + col) <= 28922) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 28923 && (row * 640 + col) <= 29281) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 29282 && (row * 640 + col) <= 29395) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 29396 && (row * 640 + col) <= 29439) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 29440 && (row * 640 + col) <= 29561) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 29562 && (row * 640 + col) <= 29923) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 29924 && (row * 640 + col) <= 30035) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 30036 && (row * 640 + col) <= 30079) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 30080 && (row * 640 + col) <= 30201) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 30202 && (row * 640 + col) <= 30562) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 30563 && (row * 640 + col) <= 30674) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 30675 && (row * 640 + col) <= 30719) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 30720 && (row * 640 + col) <= 30840) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 30841 && (row * 640 + col) <= 31202) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 31203 && (row * 640 + col) <= 31312) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31313 && (row * 640 + col) <= 31359) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 31360 && (row * 640 + col) <= 31480) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 31481 && (row * 640 + col) <= 31842) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 31843 && (row * 640 + col) <= 31951) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 31952 && (row * 640 + col) <= 31999) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 32000 && (row * 640 + col) <= 32119) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 32120 && (row * 640 + col) <= 32482) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 32483 && (row * 640 + col) <= 32589) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 32590 && (row * 640 + col) <= 32639) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 32640 && (row * 640 + col) <= 32759) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 32760 && (row * 640 + col) <= 33122) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 33123 && (row * 640 + col) <= 33226) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33227 && (row * 640 + col) <= 33279) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 33280 && (row * 640 + col) <= 33398) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 33399 && (row * 640 + col) <= 33762) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 33763 && (row * 640 + col) <= 33862) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 33863 && (row * 640 + col) <= 33919) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 33920 && (row * 640 + col) <= 34038) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 34039 && (row * 640 + col) <= 34402) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 34403 && (row * 640 + col) <= 34501) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 34502 && (row * 640 + col) <= 34559) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 34560 && (row * 640 + col) <= 34677) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 34678 && (row * 640 + col) <= 35043) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 35044 && (row * 640 + col) <= 35141) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35142 && (row * 640 + col) <= 35199) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 35200 && (row * 640 + col) <= 35317) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 35318 && (row * 640 + col) <= 35684) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 35685 && (row * 640 + col) <= 35780) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 35781 && (row * 640 + col) <= 35839) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 35840 && (row * 640 + col) <= 35956) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 35957 && (row * 640 + col) <= 36325) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 36326 && (row * 640 + col) <= 36419) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 36420 && (row * 640 + col) <= 36479) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 36480 && (row * 640 + col) <= 36596) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 36597 && (row * 640 + col) <= 36967) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 36968 && (row * 640 + col) <= 37058) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37059 && (row * 640 + col) <= 37119) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 37120 && (row * 640 + col) <= 37235) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 37236 && (row * 640 + col) <= 37609) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 37610 && (row * 640 + col) <= 37697) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 37698 && (row * 640 + col) <= 37759) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 37760 && (row * 640 + col) <= 37874) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 37875 && (row * 640 + col) <= 38253) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 38254 && (row * 640 + col) <= 38335) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38336 && (row * 640 + col) <= 38399) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 38400 && (row * 640 + col) <= 38514) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 38515 && (row * 640 + col) <= 38895) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 38896 && (row * 640 + col) <= 38972) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 38973 && (row * 640 + col) <= 39039) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 39040 && (row * 640 + col) <= 39153) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 39154 && (row * 640 + col) <= 39536) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 39537 && (row * 640 + col) <= 39598) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39599 && (row * 640 + col) <= 39602) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 39603 && (row * 640 + col) <= 39607) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 39608 && (row * 640 + col) <= 39679) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 39680 && (row * 640 + col) <= 39793) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 39794 && (row * 640 + col) <= 40182) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 40183 && (row * 640 + col) <= 40237) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40238 && (row * 640 + col) <= 40319) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 40320 && (row * 640 + col) <= 40432) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 40433 && (row * 640 + col) <= 40827) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 40828 && (row * 640 + col) <= 40843) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40844 && (row * 640 + col) <= 40844) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 40845 && (row * 640 + col) <= 40876) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 40877 && (row * 640 + col) <= 40959) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 40960 && (row * 640 + col) <= 41071) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 41072 && (row * 640 + col) <= 41469) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 41470 && (row * 640 + col) <= 41479) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 41480 && (row * 640 + col) <= 41485) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 41486 && (row * 640 + col) <= 41514) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 41515 && (row * 640 + col) <= 41599) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 41600 && (row * 640 + col) <= 41711) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 41712 && (row * 640 + col) <= 42127) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 42128 && (row * 640 + col) <= 42152) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42153 && (row * 640 + col) <= 42239) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 42240 && (row * 640 + col) <= 42350) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 42351 && (row * 640 + col) <= 42770) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 42771 && (row * 640 + col) <= 42790) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 42791 && (row * 640 + col) <= 42879) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 42880 && (row * 640 + col) <= 42989) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 42990 && (row * 640 + col) <= 43414) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 43415 && (row * 640 + col) <= 43426) color_data <= 12'b111111111111; else
        if ((row * 640 + col) >= 43427 && (row * 640 + col) <= 43519) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 43520 && (row * 640 + col) <= 43629) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 43630 && (row * 640 + col) <= 44159) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 44160 && (row * 640 + col) <= 44268) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 44269 && (row * 640 + col) <= 44799) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 44800 && (row * 640 + col) <= 44907) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 44908 && (row * 640 + col) <= 45439) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 45440 && (row * 640 + col) <= 45546) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 45547 && (row * 640 + col) <= 46079) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 46080 && (row * 640 + col) <= 46185) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 46186 && (row * 640 + col) <= 46719) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 46720 && (row * 640 + col) <= 46825) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 46826 && (row * 640 + col) <= 47359) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 47360 && (row * 640 + col) <= 47464) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 47465 && (row * 640 + col) <= 47999) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 48000 && (row * 640 + col) <= 48103) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 48104 && (row * 640 + col) <= 48639) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 48640 && (row * 640 + col) <= 48742) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 48743 && (row * 640 + col) <= 49279) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 49280 && (row * 640 + col) <= 49381) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 49382 && (row * 640 + col) <= 49919) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 49920 && (row * 640 + col) <= 50020) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 50021 && (row * 640 + col) <= 50559) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 50560 && (row * 640 + col) <= 50659) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 50660 && (row * 640 + col) <= 51199) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 51200 && (row * 640 + col) <= 51298) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 51299 && (row * 640 + col) <= 51839) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 51840 && (row * 640 + col) <= 51937) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 51938 && (row * 640 + col) <= 52479) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 52480 && (row * 640 + col) <= 52576) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 52577 && (row * 640 + col) <= 53119) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 53120 && (row * 640 + col) <= 53215) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 53216 && (row * 640 + col) <= 53759) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 53760 && (row * 640 + col) <= 53854) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 53855 && (row * 640 + col) <= 54399) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 54400 && (row * 640 + col) <= 54493) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 54494 && (row * 640 + col) <= 55039) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 55040 && (row * 640 + col) <= 55132) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 55133 && (row * 640 + col) <= 55679) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 55680 && (row * 640 + col) <= 55771) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 55772 && (row * 640 + col) <= 56319) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 56320 && (row * 640 + col) <= 56410) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 56411 && (row * 640 + col) <= 56959) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 56960 && (row * 640 + col) <= 57049) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 57050 && (row * 640 + col) <= 57599) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 57600 && (row * 640 + col) <= 57688) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 57689 && (row * 640 + col) <= 58239) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 58240 && (row * 640 + col) <= 58326) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 58327 && (row * 640 + col) <= 58879) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 58880 && (row * 640 + col) <= 58965) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 58966 && (row * 640 + col) <= 59519) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 59520 && (row * 640 + col) <= 59604) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 59605 && (row * 640 + col) <= 60159) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 60160 && (row * 640 + col) <= 60243) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 60244 && (row * 640 + col) <= 60799) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 60800 && (row * 640 + col) <= 60881) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 60882 && (row * 640 + col) <= 61439) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 61440 && (row * 640 + col) <= 61520) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 61521 && (row * 640 + col) <= 62079) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 62080 && (row * 640 + col) <= 62158) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 62159 && (row * 640 + col) <= 62719) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 62720 && (row * 640 + col) <= 62797) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 62798 && (row * 640 + col) <= 63359) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 63360 && (row * 640 + col) <= 63436) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 63437 && (row * 640 + col) <= 63999) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 64000 && (row * 640 + col) <= 64074) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 64075 && (row * 640 + col) <= 64639) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 64640 && (row * 640 + col) <= 64713) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 64714 && (row * 640 + col) <= 65279) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 65280 && (row * 640 + col) <= 65351) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 65352 && (row * 640 + col) <= 65919) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 65920 && (row * 640 + col) <= 65989) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 65990 && (row * 640 + col) <= 66559) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 66560 && (row * 640 + col) <= 66627) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 66628 && (row * 640 + col) <= 67199) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 67200 && (row * 640 + col) <= 67265) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 67266 && (row * 640 + col) <= 67839) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 67840 && (row * 640 + col) <= 67904) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 67905 && (row * 640 + col) <= 68479) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 68480 && (row * 640 + col) <= 68542) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 68543 && (row * 640 + col) <= 69119) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 69120 && (row * 640 + col) <= 69180) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 69181 && (row * 640 + col) <= 69759) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 69760 && (row * 640 + col) <= 69817) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 69818 && (row * 640 + col) <= 70399) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 70400 && (row * 640 + col) <= 70455) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 70456 && (row * 640 + col) <= 71039) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 71040 && (row * 640 + col) <= 71093) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 71094 && (row * 640 + col) <= 71679) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 71680 && (row * 640 + col) <= 71731) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 71732 && (row * 640 + col) <= 72319) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 72320 && (row * 640 + col) <= 72368) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 72369 && (row * 640 + col) <= 72959) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 72960 && (row * 640 + col) <= 73005) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 73006 && (row * 640 + col) <= 73599) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 73600 && (row * 640 + col) <= 73642) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 73643 && (row * 640 + col) <= 74239) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 74240 && (row * 640 + col) <= 74279) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 74280 && (row * 640 + col) <= 74879) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 74880 && (row * 640 + col) <= 74914) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 74915 && (row * 640 + col) <= 75519) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 75520 && (row * 640 + col) <= 75550) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 75551 && (row * 640 + col) <= 76159) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 76160 && (row * 640 + col) <= 76186) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 76187 && (row * 640 + col) <= 76799) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 76800 && (row * 640 + col) <= 76819) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 76820 && (row * 640 + col) <= 77439) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 77440 && (row * 640 + col) <= 77450) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 77451 && (row * 640 + col) <= 202879) color_data <= 12'b000010101110; else
        if ((row * 640 + col) >= 202880 && (row * 640 + col) <= 226559) color_data <= 12'b001010110100; else
        if ((row * 640 + col) >= 226560 && (row * 640 + col) <= 249364) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249365 && (row * 640 + col) <= 249407) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 249408 && (row * 640 + col) <= 249515) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249516 && (row * 640 + col) <= 249558) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 249559 && (row * 640 + col) <= 249927) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 249928 && (row * 640 + col) <= 249970) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 249971 && (row * 640 + col) <= 250004) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250005 && (row * 640 + col) <= 250047) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250048 && (row * 640 + col) <= 250083) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250084 && (row * 640 + col) <= 250126) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250127 && (row * 640 + col) <= 250155) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250156 && (row * 640 + col) <= 250198) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250199 && (row * 640 + col) <= 250266) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250267 && (row * 640 + col) <= 250309) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250310 && (row * 640 + col) <= 250337) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250338 && (row * 640 + col) <= 250380) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250381 && (row * 640 + col) <= 250485) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250486 && (row * 640 + col) <= 250528) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250529 && (row * 640 + col) <= 250567) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250568 && (row * 640 + col) <= 250610) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250611 && (row * 640 + col) <= 250644) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250645 && (row * 640 + col) <= 250687) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250688 && (row * 640 + col) <= 250723) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250724 && (row * 640 + col) <= 250766) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250767 && (row * 640 + col) <= 250795) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250796 && (row * 640 + col) <= 250838) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250839 && (row * 640 + col) <= 250906) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250907 && (row * 640 + col) <= 250949) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 250950 && (row * 640 + col) <= 250977) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 250978 && (row * 640 + col) <= 251020) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251021 && (row * 640 + col) <= 251050) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251051 && (row * 640 + col) <= 251093) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251094 && (row * 640 + col) <= 251125) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251126 && (row * 640 + col) <= 251168) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251169 && (row * 640 + col) <= 251207) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251208 && (row * 640 + col) <= 251250) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251251 && (row * 640 + col) <= 251284) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251285 && (row * 640 + col) <= 251327) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251328 && (row * 640 + col) <= 251363) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251364 && (row * 640 + col) <= 251406) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251407 && (row * 640 + col) <= 251435) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251436 && (row * 640 + col) <= 251478) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251479 && (row * 640 + col) <= 251546) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251547 && (row * 640 + col) <= 251589) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251590 && (row * 640 + col) <= 251617) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251618 && (row * 640 + col) <= 251660) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251661 && (row * 640 + col) <= 251690) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251691 && (row * 640 + col) <= 251733) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251734 && (row * 640 + col) <= 251765) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251766 && (row * 640 + col) <= 251808) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251809 && (row * 640 + col) <= 251847) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251848 && (row * 640 + col) <= 251890) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251891 && (row * 640 + col) <= 251924) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 251925 && (row * 640 + col) <= 251967) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 251968 && (row * 640 + col) <= 252003) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252004 && (row * 640 + col) <= 252046) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252047 && (row * 640 + col) <= 252075) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252076 && (row * 640 + col) <= 252118) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252119 && (row * 640 + col) <= 252186) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252187 && (row * 640 + col) <= 252229) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252230 && (row * 640 + col) <= 252257) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252258 && (row * 640 + col) <= 252300) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252301 && (row * 640 + col) <= 252330) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252331 && (row * 640 + col) <= 252373) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252374 && (row * 640 + col) <= 252405) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252406 && (row * 640 + col) <= 252448) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252449 && (row * 640 + col) <= 252487) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252488 && (row * 640 + col) <= 252530) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252531 && (row * 640 + col) <= 252564) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252565 && (row * 640 + col) <= 252607) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252608 && (row * 640 + col) <= 252643) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252644 && (row * 640 + col) <= 252686) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252687 && (row * 640 + col) <= 252715) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252716 && (row * 640 + col) <= 252758) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252759 && (row * 640 + col) <= 252826) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252827 && (row * 640 + col) <= 252869) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252870 && (row * 640 + col) <= 252897) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252898 && (row * 640 + col) <= 252940) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 252941 && (row * 640 + col) <= 252970) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 252971 && (row * 640 + col) <= 253013) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253014 && (row * 640 + col) <= 253045) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253046 && (row * 640 + col) <= 253088) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253089 && (row * 640 + col) <= 253127) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253128 && (row * 640 + col) <= 253170) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253171 && (row * 640 + col) <= 253204) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253205 && (row * 640 + col) <= 253247) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253248 && (row * 640 + col) <= 253283) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253284 && (row * 640 + col) <= 253326) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253327 && (row * 640 + col) <= 253355) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253356 && (row * 640 + col) <= 253398) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253399 && (row * 640 + col) <= 253466) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253467 && (row * 640 + col) <= 253509) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253510 && (row * 640 + col) <= 253537) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253538 && (row * 640 + col) <= 253580) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253581 && (row * 640 + col) <= 253610) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253611 && (row * 640 + col) <= 253653) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253654 && (row * 640 + col) <= 253685) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253686 && (row * 640 + col) <= 253728) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253729 && (row * 640 + col) <= 253767) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253768 && (row * 640 + col) <= 253810) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253811 && (row * 640 + col) <= 253844) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253845 && (row * 640 + col) <= 253887) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253888 && (row * 640 + col) <= 253923) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253924 && (row * 640 + col) <= 253966) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 253967 && (row * 640 + col) <= 253995) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 253996 && (row * 640 + col) <= 254038) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254039 && (row * 640 + col) <= 254106) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254107 && (row * 640 + col) <= 254149) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254150 && (row * 640 + col) <= 254177) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254178 && (row * 640 + col) <= 254220) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254221 && (row * 640 + col) <= 254250) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254251 && (row * 640 + col) <= 254293) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254294 && (row * 640 + col) <= 254325) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254326 && (row * 640 + col) <= 254368) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254369 && (row * 640 + col) <= 254407) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254408 && (row * 640 + col) <= 254450) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254451 && (row * 640 + col) <= 254484) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254485 && (row * 640 + col) <= 254527) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254528 && (row * 640 + col) <= 254563) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254564 && (row * 640 + col) <= 254606) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254607 && (row * 640 + col) <= 254635) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254636 && (row * 640 + col) <= 254678) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254679 && (row * 640 + col) <= 254746) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254747 && (row * 640 + col) <= 254789) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254790 && (row * 640 + col) <= 254817) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254818 && (row * 640 + col) <= 254860) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254861 && (row * 640 + col) <= 254890) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254891 && (row * 640 + col) <= 254933) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 254934 && (row * 640 + col) <= 254965) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 254966 && (row * 640 + col) <= 255008) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255009 && (row * 640 + col) <= 255047) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255048 && (row * 640 + col) <= 255090) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255091 && (row * 640 + col) <= 255124) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255125 && (row * 640 + col) <= 255167) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255168 && (row * 640 + col) <= 255203) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255204 && (row * 640 + col) <= 255246) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255247 && (row * 640 + col) <= 255275) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255276 && (row * 640 + col) <= 255318) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255319 && (row * 640 + col) <= 255386) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255387 && (row * 640 + col) <= 255429) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255430 && (row * 640 + col) <= 255457) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255458 && (row * 640 + col) <= 255500) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255501 && (row * 640 + col) <= 255530) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255531 && (row * 640 + col) <= 255573) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255574 && (row * 640 + col) <= 255605) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255606 && (row * 640 + col) <= 255648) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255649 && (row * 640 + col) <= 255687) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255688 && (row * 640 + col) <= 255730) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255731 && (row * 640 + col) <= 255764) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255765 && (row * 640 + col) <= 255807) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255808 && (row * 640 + col) <= 255843) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255844 && (row * 640 + col) <= 255886) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255887 && (row * 640 + col) <= 255915) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 255916 && (row * 640 + col) <= 255958) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 255959 && (row * 640 + col) <= 256026) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256027 && (row * 640 + col) <= 256069) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256070 && (row * 640 + col) <= 256097) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256098 && (row * 640 + col) <= 256140) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256141 && (row * 640 + col) <= 256170) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256171 && (row * 640 + col) <= 256213) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256214 && (row * 640 + col) <= 256245) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256246 && (row * 640 + col) <= 256288) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256289 && (row * 640 + col) <= 256327) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256328 && (row * 640 + col) <= 256370) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256371 && (row * 640 + col) <= 256483) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256484 && (row * 640 + col) <= 256526) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256527 && (row * 640 + col) <= 256666) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256667 && (row * 640 + col) <= 256709) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256710 && (row * 640 + col) <= 256737) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256738 && (row * 640 + col) <= 256780) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256781 && (row * 640 + col) <= 256810) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256811 && (row * 640 + col) <= 256853) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256854 && (row * 640 + col) <= 256885) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 256886 && (row * 640 + col) <= 256928) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 256929 && (row * 640 + col) <= 257450) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 257451 && (row * 640 + col) <= 257493) color_data <= 12'b111111110000; else
        if ((row * 640 + col) >= 257494 && (row * 640 + col) <= 279679) color_data <= 12'b000000000000; else
        if ((row * 640 + col) >= 279680 && (row * 640 + col) < 307200) color_data <= 12'b001010110100; else
        color_data <= 12'b000000000000;
    end
endmodule
