module dead_player_rom (
	input wire clk,
    input wire [6:0] row,
    input wire [6:0] col,
    output reg [11:0] color_data
);

    always @(posedge clk) begin
        if ((row * 92 + col) >= 0 && (row * 92 + col) <= 117) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 125 && (row * 92 + col) <= 209) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 211 && (row * 92 + col) <= 215) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 217 && (row * 92 + col) <= 301) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 303 && (row * 92 + col) <= 307) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 309 && (row * 92 + col) <= 393) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 395 && (row * 92 + col) <= 399) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 401 && (row * 92 + col) <= 485) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 487 && (row * 92 + col) <= 491) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 493 && (row * 92 + col) <= 577) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 579 && (row * 92 + col) <= 583) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 585 && (row * 92 + col) <= 669) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 671 && (row * 92 + col) <= 675) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 677 && (row * 92 + col) <= 761) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 763 && (row * 92 + col) <= 767) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 769 && (row * 92 + col) <= 853) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 855 && (row * 92 + col) <= 859) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 861 && (row * 92 + col) <= 945) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 947 && (row * 92 + col) <= 951) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 953 && (row * 92 + col) <= 1037) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1039 && (row * 92 + col) <= 1043) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1045 && (row * 92 + col) <= 1129) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1131 && (row * 92 + col) <= 1135) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1137 && (row * 92 + col) <= 1221) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1223 && (row * 92 + col) <= 1227) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1229 && (row * 92 + col) <= 1313) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1315 && (row * 92 + col) <= 1319) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1321 && (row * 92 + col) <= 1405) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1407 && (row * 92 + col) <= 1411) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1413 && (row * 92 + col) <= 1497) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1499 && (row * 92 + col) <= 1503) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1505 && (row * 92 + col) <= 1589) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1591 && (row * 92 + col) <= 1595) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1597 && (row * 92 + col) <= 1646) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1655 && (row * 92 + col) <= 1681) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1683 && (row * 92 + col) <= 1687) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1689 && (row * 92 + col) <= 1738) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1740 && (row * 92 + col) <= 1745) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 1747 && (row * 92 + col) <= 1773) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1775 && (row * 92 + col) <= 1779) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1781 && (row * 92 + col) <= 1830) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1832 && (row * 92 + col) <= 1837) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 1839 && (row * 92 + col) <= 1865) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1867 && (row * 92 + col) <= 1871) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1873 && (row * 92 + col) <= 1922) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1924 && (row * 92 + col) <= 1929) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 1931 && (row * 92 + col) <= 1957) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 1959 && (row * 92 + col) <= 1963) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 1965 && (row * 92 + col) <= 2014) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2016 && (row * 92 + col) <= 2021) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2023 && (row * 92 + col) <= 2049) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2051 && (row * 92 + col) <= 2055) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 2057 && (row * 92 + col) <= 2106) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2108 && (row * 92 + col) <= 2113) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2115 && (row * 92 + col) <= 2141) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2143 && (row * 92 + col) <= 2147) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2149 && (row * 92 + col) <= 2198) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2200 && (row * 92 + col) <= 2205) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2207 && (row * 92 + col) <= 2233) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2235 && (row * 92 + col) <= 2239) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2241 && (row * 92 + col) <= 2290) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2292 && (row * 92 + col) <= 2297) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2299 && (row * 92 + col) <= 2325) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2327 && (row * 92 + col) <= 2331) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2333 && (row * 92 + col) <= 2382) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2384 && (row * 92 + col) <= 2389) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2391 && (row * 92 + col) <= 2417) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2419 && (row * 92 + col) <= 2423) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2425 && (row * 92 + col) <= 2474) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2476 && (row * 92 + col) <= 2481) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2483 && (row * 92 + col) <= 2509) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2511 && (row * 92 + col) <= 2515) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2517 && (row * 92 + col) <= 2566) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2568 && (row * 92 + col) <= 2573) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2575 && (row * 92 + col) <= 2601) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2603 && (row * 92 + col) <= 2607) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2660 && (row * 92 + col) <= 2665) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2667 && (row * 92 + col) <= 2678) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2685 && (row * 92 + col) <= 2693) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2695 && (row * 92 + col) <= 2728) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2729 && (row * 92 + col) <= 2750) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 2751 && (row * 92 + col) <= 2757) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2759 && (row * 92 + col) <= 2766) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2771 && (row * 92 + col) <= 2776) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 2780 && (row * 92 + col) <= 2785) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2787 && (row * 92 + col) <= 2820) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2821 && (row * 92 + col) <= 2842) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 2843 && (row * 92 + col) <= 2849) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2851 && (row * 92 + col) <= 2858) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2860 && (row * 92 + col) <= 2871) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 2873 && (row * 92 + col) <= 2877) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2879 && (row * 92 + col) <= 2912) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 2913 && (row * 92 + col) <= 2934) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 2935 && (row * 92 + col) <= 2941) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 2943 && (row * 92 + col) <= 2948) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2951 && (row * 92 + col) <= 2964) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 2967 && (row * 92 + col) <= 2969) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 2971 && (row * 92 + col) <= 3004) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3005 && (row * 92 + col) <= 3026) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3027 && (row * 92 + col) <= 3033) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 3035 && (row * 92 + col) <= 3039) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3041 && (row * 92 + col) <= 3058) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3060 && (row * 92 + col) <= 3061) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3063 && (row * 92 + col) <= 3096) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3097 && (row * 92 + col) <= 3118) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3119 && (row * 92 + col) <= 3125) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 3127 && (row * 92 + col) <= 3131) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3133 && (row * 92 + col) <= 3150) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3152 && (row * 92 + col) <= 3153) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3155 && (row * 92 + col) <= 3188) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3189 && (row * 92 + col) <= 3210) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3211 && (row * 92 + col) <= 3217) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 3219 && (row * 92 + col) <= 3222) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3224 && (row * 92 + col) <= 3243) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3245 && (row * 92 + col) <= 3245) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3247 && (row * 92 + col) <= 3280) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3281 && (row * 92 + col) <= 3285) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3311 && (row * 92 + col) <= 3313) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3315 && (row * 92 + col) <= 3318) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3320 && (row * 92 + col) <= 3322) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3324 && (row * 92 + col) <= 3331) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3334 && (row * 92 + col) <= 3336) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3339 && (row * 92 + col) <= 3372) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3373 && (row * 92 + col) <= 3377) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3379 && (row * 92 + col) <= 3405) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3407 && (row * 92 + col) <= 3411) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3413 && (row * 92 + col) <= 3413) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3415 && (row * 92 + col) <= 3422) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3426 && (row * 92 + col) <= 3429) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3431 && (row * 92 + col) <= 3464) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3465 && (row * 92 + col) <= 3469) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3471 && (row * 92 + col) <= 3497) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3499 && (row * 92 + col) <= 3504) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3506 && (row * 92 + col) <= 3513) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3516 && (row * 92 + col) <= 3516) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 3518 && (row * 92 + col) <= 3522) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3523 && (row * 92 + col) <= 3556) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3557 && (row * 92 + col) <= 3561) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3563 && (row * 92 + col) <= 3588) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3590 && (row * 92 + col) <= 3595) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3597 && (row * 92 + col) <= 3597) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3599 && (row * 92 + col) <= 3605) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3607 && (row * 92 + col) <= 3608) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 3610 && (row * 92 + col) <= 3614) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3615 && (row * 92 + col) <= 3648) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3649 && (row * 92 + col) <= 3653) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3655 && (row * 92 + col) <= 3680) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3682 && (row * 92 + col) <= 3686) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3688 && (row * 92 + col) <= 3690) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3692 && (row * 92 + col) <= 3697) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3699 && (row * 92 + col) <= 3700) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 3702 && (row * 92 + col) <= 3706) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3707 && (row * 92 + col) <= 3740) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3741 && (row * 92 + col) <= 3745) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3747 && (row * 92 + col) <= 3772) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3774 && (row * 92 + col) <= 3788) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3791 && (row * 92 + col) <= 3792) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 3794 && (row * 92 + col) <= 3798) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3799 && (row * 92 + col) <= 3832) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3833 && (row * 92 + col) <= 3837) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3839 && (row * 92 + col) <= 3864) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3866 && (row * 92 + col) <= 3880) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3882 && (row * 92 + col) <= 3884) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 3886 && (row * 92 + col) <= 3890) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3891 && (row * 92 + col) <= 3924) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 3925 && (row * 92 + col) <= 3929) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 3931 && (row * 92 + col) <= 3956) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 3958 && (row * 92 + col) <= 3972) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3974 && (row * 92 + col) <= 3976) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 3978 && (row * 92 + col) <= 3982) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 3983 && (row * 92 + col) <= 4016) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4017 && (row * 92 + col) <= 4021) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4023 && (row * 92 + col) <= 4048) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4050 && (row * 92 + col) <= 4054) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4056 && (row * 92 + col) <= 4058) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4060 && (row * 92 + col) <= 4064) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4066 && (row * 92 + col) <= 4068) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 4070 && (row * 92 + col) <= 4074) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4075 && (row * 92 + col) <= 4108) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4109 && (row * 92 + col) <= 4113) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4115 && (row * 92 + col) <= 4141) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4143 && (row * 92 + col) <= 4147) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4149 && (row * 92 + col) <= 4149) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4151 && (row * 92 + col) <= 4156) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4159 && (row * 92 + col) <= 4160) color_data <= 12'b111011101110; else
        if ((row * 92 + col) >= 4162 && (row * 92 + col) <= 4166) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4167 && (row * 92 + col) <= 4200) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4201 && (row * 92 + col) <= 4205) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4207 && (row * 92 + col) <= 4233) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4235 && (row * 92 + col) <= 4240) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4242 && (row * 92 + col) <= 4249) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4254 && (row * 92 + col) <= 4257) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4259 && (row * 92 + col) <= 4292) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4293 && (row * 92 + col) <= 4297) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4323 && (row * 92 + col) <= 4325) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4327 && (row * 92 + col) <= 4331) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4333 && (row * 92 + col) <= 4333) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4335 && (row * 92 + col) <= 4343) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4346 && (row * 92 + col) <= 4348) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4351 && (row * 92 + col) <= 4384) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4385 && (row * 92 + col) <= 4406) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4407 && (row * 92 + col) <= 4413) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 4415 && (row * 92 + col) <= 4418) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4420 && (row * 92 + col) <= 4422) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4424 && (row * 92 + col) <= 4426) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4428 && (row * 92 + col) <= 4439) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4441 && (row * 92 + col) <= 4441) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4443 && (row * 92 + col) <= 4476) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4477 && (row * 92 + col) <= 4498) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4499 && (row * 92 + col) <= 4505) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 4507 && (row * 92 + col) <= 4511) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4513 && (row * 92 + col) <= 4530) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4532 && (row * 92 + col) <= 4533) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4535 && (row * 92 + col) <= 4568) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4569 && (row * 92 + col) <= 4590) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4591 && (row * 92 + col) <= 4597) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 4599 && (row * 92 + col) <= 4603) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4605 && (row * 92 + col) <= 4622) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4624 && (row * 92 + col) <= 4625) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4627 && (row * 92 + col) <= 4660) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4661 && (row * 92 + col) <= 4682) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4683 && (row * 92 + col) <= 4689) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 4691 && (row * 92 + col) <= 4696) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4699 && (row * 92 + col) <= 4712) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4715 && (row * 92 + col) <= 4717) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4719 && (row * 92 + col) <= 4752) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4753 && (row * 92 + col) <= 4774) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4775 && (row * 92 + col) <= 4781) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 4783 && (row * 92 + col) <= 4790) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4793 && (row * 92 + col) <= 4803) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4805 && (row * 92 + col) <= 4809) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4811 && (row * 92 + col) <= 4844) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4845 && (row * 92 + col) <= 4866) color_data <= 12'b001101001100; else
        if ((row * 92 + col) >= 4867 && (row * 92 + col) <= 4873) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 4875 && (row * 92 + col) <= 4884) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4887 && (row * 92 + col) <= 4892) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 4896 && (row * 92 + col) <= 4901) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4903 && (row * 92 + col) <= 4907) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 4960 && (row * 92 + col) <= 4965) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 4967 && (row * 92 + col) <= 4978) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4985 && (row * 92 + col) <= 4993) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 4995 && (row * 92 + col) <= 4999) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 5001 && (row * 92 + col) <= 5050) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5052 && (row * 92 + col) <= 5057) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5059 && (row * 92 + col) <= 5085) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5087 && (row * 92 + col) <= 5091) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 5093 && (row * 92 + col) <= 5142) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5144 && (row * 92 + col) <= 5149) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5151 && (row * 92 + col) <= 5177) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5179 && (row * 92 + col) <= 5183) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 5185 && (row * 92 + col) <= 5234) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5236 && (row * 92 + col) <= 5241) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5243 && (row * 92 + col) <= 5269) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5271 && (row * 92 + col) <= 5275) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 5277 && (row * 92 + col) <= 5326) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5328 && (row * 92 + col) <= 5333) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5335 && (row * 92 + col) <= 5361) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5363 && (row * 92 + col) <= 5367) color_data <= 12'b111000010010; else
        if ((row * 92 + col) >= 5369 && (row * 92 + col) <= 5418) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5420 && (row * 92 + col) <= 5425) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5427 && (row * 92 + col) <= 5453) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5455 && (row * 92 + col) <= 5459) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 5461 && (row * 92 + col) <= 5510) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5512 && (row * 92 + col) <= 5517) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5519 && (row * 92 + col) <= 5545) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5547 && (row * 92 + col) <= 5551) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 5553 && (row * 92 + col) <= 5602) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5604 && (row * 92 + col) <= 5609) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5611 && (row * 92 + col) <= 5637) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5639 && (row * 92 + col) <= 5643) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 5645 && (row * 92 + col) <= 5694) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5696 && (row * 92 + col) <= 5701) color_data <= 12'b101101110101; else
        if ((row * 92 + col) >= 5703 && (row * 92 + col) <= 5729) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5731 && (row * 92 + col) <= 5735) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 5737 && (row * 92 + col) <= 5786) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5795 && (row * 92 + col) <= 5821) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5823 && (row * 92 + col) <= 5827) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 5829 && (row * 92 + col) <= 5913) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 5915 && (row * 92 + col) <= 5919) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 5921 && (row * 92 + col) <= 6005) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6007 && (row * 92 + col) <= 6011) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6013 && (row * 92 + col) <= 6097) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6099 && (row * 92 + col) <= 6103) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6105 && (row * 92 + col) <= 6189) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6191 && (row * 92 + col) <= 6195) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6197 && (row * 92 + col) <= 6281) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6283 && (row * 92 + col) <= 6287) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6289 && (row * 92 + col) <= 6373) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6375 && (row * 92 + col) <= 6379) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6381 && (row * 92 + col) <= 6465) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6467 && (row * 92 + col) <= 6471) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6473 && (row * 92 + col) <= 6557) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6559 && (row * 92 + col) <= 6563) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6565 && (row * 92 + col) <= 6649) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6651 && (row * 92 + col) <= 6655) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6657 && (row * 92 + col) <= 6741) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6743 && (row * 92 + col) <= 6747) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6749 && (row * 92 + col) <= 6833) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6835 && (row * 92 + col) <= 6839) color_data <= 12'b111111111010; else
        if ((row * 92 + col) >= 6841 && (row * 92 + col) <= 6925) color_data <= 12'b111111111111; else
        if ((row * 92 + col) >= 6933 && (row * 92 + col) < 7084) color_data <= 12'b111111111111; else
        color_data <= 12'b000000000000;
    end
endmodule